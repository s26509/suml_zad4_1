���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.6.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy._core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h3�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh'�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M�nodes�h)h,K ��h.��R�(KM��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h~h3�i8�����R�(KhMNNNJ����J����K t�bK ��hh�K��h�h�K��h�h^K��h�h^K ��h�h�K(��h�h^K0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@E         �                     @"��p�?�           8�@               u                    �?.y0��k�?�            �s@              "                    �?Hث3���?�            @m@                                   �?     ��?)             P@                               0�FF@�'N��?&            �N@                                 s�,@�q�����?             9@        ������������������������       �                     @               	                 �܅3@8�A�0��?             6@        ������������������������       �                     @        
                        p�i@@�\��N��?             3@                                  �?��
ц��?	             *@                                   �?      �?             @        ������������������������       �                     �?                                  �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �<@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                                   �?�����H�?             B@       ������������������������       �                     9@                                p"�X@���|���?             &@                                 �8@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                !                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        #       &                   �9@���Q��?i            @e@        $       %                    �?��s����?             5@        ������������������������       �                     @        ������������������������       �                     1@        '       f                  x#J@p�B<F]�?[            �b@       (       G                     �?��c`��?L            �^@        )       >                   �>@8����?              G@       *       +                    �?��
ц��?             :@        ������������������������       �                     @        ,       -                   �<@�q�q�?             5@        ������������������������       �                     @        .       =                    R@�<ݚ�?             2@       /       0                 03:@@�0�!��?             1@        ������������������������       �                     @        1       <                   �J@���!pc�?	             &@       2       3                 03k:@      �?              @        ������������������������       �                     �?        4       ;                    H@����X�?             @       5       :                 X��B@r�q��?             @       6       7                 `fF<@      �?             @        ������������������������       �                      @        8       9                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ?       @                 `f~I@ףp=
�?             4@       ������������������������       �                     (@        A       B                 `��I@      �?              @        ������������������������       �                     �?        C       D                 03�I@؇���X�?             @        ������������������������       �                     �?        E       F                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        H       e                    >@&:~�Q�?,             S@       I       X                    �?�Y�R_�?+            �Q@        J       K                   @B@ �o_��?             9@        ������������������������       �                     "@        L       S                    -@     ��?             0@       M       P                   �'@      �?              @        N       O                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Q       R                    D@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        T       W                   �H@      �?              @       U       V                   �E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Y       d                    �?���}<S�?             G@       Z       c                   @A@��-�=��?            �C@        [       b                   �@@������?
             1@       \       ]                 �|Y=@�r����?	             .@        ������������������������       �                     @        ^       _                   �'@�<ݚ�?             "@       ������������������������       �                     @        `       a                 �|�=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     @        ������������������������       �                     @        g       t                 03�U@PN��T'�?             ;@       h       i                    <@��s����?             5@        ������������������������       �                     @        j       k                    ?@      �?	             0@        ������������������������       �                     �?        l       m                    B@z�G�z�?             .@        ������������������������       �                     @        n       o                    C@�z�G��?             $@        ������������������������       �                      @        p       q                    �?      �?              @        ������������������������       �                     @        r       s                 0� Q@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    :@���B���?3            �S@        ������������������������       �        
             1@        x                          �8@�jTM��?)            �N@        y       ~                    @�g�y��?             ?@        z       {                 ��W@      �?             @        ������������������������       �                      @        |       }                 �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    �?��S���?             >@       �       �                  DT@�ՙ/�?             5@       �       �                     �?�n_Y�K�?	             *@        �       �                 X�,D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �UA@r�q��?             @       �       �                   @A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�~�@
�?�            �x@        �       �                    7@�g�y��?             ?@        �       �                 03�@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     5@        �       
                ��Y7@�?��+�?�             w@       �       �                    /@����I�?�            �t@        �       �                    $@      �?             8@       ������������������������       �        	             .@        �       �                 �&�)@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����Y��?�            s@        �       �                    �?���ȫ�?/            �T@        �       �                    �?�MI8d�?            �B@       �       �                    �?      �?             @@       ������������������������       �                     6@        �       �                  S�-@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                 `�@1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @X�<ݚ�?            �F@       �       �                  s@~�4_�g�?             F@        ������������������������       �                     @        �       �                   �3@      �?             D@        ������������������������       �                     �?        �       �                   �4@�99lMt�?            �C@        ������������������������       �                     @        �       �                 ��/@b�2�tk�?             B@       �       �                    �?�z�G��?             >@       �       �                   �5@�û��|�?             7@        ������������������������       �                     �?        �       �                    �?���|���?             6@       �       �                   P&@�q�q�?             5@       �       �                 �|�;@�z�G��?             4@       �       �                 pf�@�n_Y�K�?             *@        ������������������������       �                      @        �       �                 pf� @���!pc�?             &@       �       �                   �9@և���X�?             @       �       �                   �6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��� @؇���X�?             @       ������������������������       �                     @        �       �                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@�@+��?�            �k@        �       �                    �?�<ݚ�?             2@       �       �                   @@$�q-�?
             *@        �       �                 �|�:@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     "@        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�M��?}            �i@        �       �                    �?XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        �       �                 �?�@h�V���?l             f@        �       �                   �?@�k~X��?.             R@       ������������������������       �        %             L@        �       �                   @@@      �?	             0@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �1@�ջ����?>             Z@        ������������������������       �                     (@        �       	                   �?��H�?7             W@       �                          �?z�G�z�?2            @U@       �       �                 @3�@*�s���?1             U@        �       �                   �?@      �?             ,@        �       �                   �9@�q�q�?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �A@      �?              @        ������������������������       ��q�q�?             @        ������������������������       ����Q��?             @        �       �                   �2@؇���X�?*            �Q@        ������������������������       �                     @        �       �                 ��) @pH����?)            �P@        �       �                   �3@ 7���B�?             ;@        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   �9@R���Q�?             D@        ������������������������       �                     1@        �                          (@��+7��?             7@       �                          ?@���Q��?             .@                              �|Y=@      �?              @        ������������������������       �                     @                              �̜!@���Q��?             @        ������������������������       �                     �?                              �|�=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                              ��T?@��-�=��?            �C@       ������������������������       �                     9@                                 �?����X�?             ,@        ������������������������       �                     @                                 @���|���?             &@                                @���Q��?             $@                             ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�b�values�h)h,K ��h.��R�(KMKK��h^�BP  J54v��?l�����?;�;��?vb'vb'�?�i�i�?��-��-�?      �?      �?ާ�d��?�����?�p=
ף�?���Q��?              �?颋.���?/�袋.�?      �?        y�5���?�5��P�?�؉�؉�?�;�;�?      �?      �?      �?        �������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?z��y���?�a�a�?              �?      �?        :��IA�?�3�=l}�?2�h�>�?��).��?d!Y�B�?8��Moz�?�;�;�?�؉�؉�?              �?UUUUUU�?UUUUUU�?              �?9��8���?�q�q�?ZZZZZZ�?�������?      �?        F]t�E�?t�E]t�?      �?      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?      �?                      �?      �?                      �?�������?�������?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?        �k(���?�k(����?���@��?�z2~���?�Q����?
ףp=
�?              �?      �?      �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?ӛ���7�?d!Y�B�?}˷|˷�?�A�A�?xxxxxx�?�?�������?�?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?                      �?h/�����?&���^B�?�a�a�?z��y���?              �?      �?      �?      �?        �������?�������?              �?333333�?ffffff�?      �?              �?      �?              �?      �?      �?              �?      �?                      �?ى�؉��?��؉���?              �?.�u�y�?�y��!�?�B!��?��{���?      �?      �?              �?      �?      �?              �?      �?                      �?�������?�?�a�a�?�<��<��?;�;��?ى�؉��?      �?      �?              �?      �?        r�q��?�q�q�?              �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?      �?              �?      �?              �?        ������?� �D
�?��{���?�B!��?�������?�������?      �?                      �?      �?        ���,d�?ӛ���7�?�|`d���??7�z�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?E�n<�?�ƃ�D�?28��1�?�cp>��?L�Ϻ��?��L���?      �?      �?              �?�������?�������?      �?                      �?�������?�������?      �?                      �?r�q��?�q�q�?/�袋.�?��.���?              �?      �?      �?              �?5H�4H��?�o��o��?      �?        �8��8��?9��8���?ffffff�?333333�?8��Moz�?��,d!�?              �?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?ffffff�?333333�?;�;��?ى�؉��?              �?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?              �?      �?        UUUUUU�?�������?      �?                      �?              �?������?;Ӹ�Qg�?9��8���?�q�q�?�؉�؉�?;�;��?      �?      �?      �?              �?      �?      �?        �������?333333�?      �?                      �?	݋н�?��{��?GX�i���?�{a���?      �?                      �?�袋.��?/�袋.�?�8��8��?�q�q�?      �?              �?      �?      �?      �?              �?      �?              �?        O��N���?�N��N��?      �?        !Y�B�?zӛ����?�������?�������?b�a��?z��y���?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?333333�?�������?۶m۶m�?�$I�$I�?              �?�1���?z�rv��?	�%����?h/�����?              �?      �?        333333�?333333�?      �?        zӛ����?Y�B��?333333�?�������?      �?      �?              �?�������?333333�?              �?      �?      �?      �?                      �?      �?              �?              �?              �?        }˷|˷�?�A�A�?      �?        �m۶m��?�$I�$I�?      �?        ]t�E]�?F]t�E�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK���h}�B�?                             @���*1�?�           8�@                                   @�7����?            �G@                                   �?Pa�	�?            �@@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@               	                 ��T?@؇���X�?             ,@        ������������������������       �                      @        
                           @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               z                     @��?a�?�           ��@               !                    �?V$�݆��?�            �r@                                 0Cd=@Pns��ޭ?O            �`@                                  @E@$Q�q�?"            �O@                               ���*@p���?             I@                                `f�)@�IєX�?	             1@        ������������������������       �                     (@                                   :@z�G�z�?             @                                   5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@                                   �?�θ�?             *@                               ���;@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        -            �Q@        "       y                    �?4>���?t             e@       #       8                 `ff:@�{��?��?n            @d@        $       '                    5@ >�֕�?0            �Q@        %       &                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                 �|Y=@ =[y��?.             Q@        ������������������������       �                     4@        *       7                   �*@      �?#             H@       +       ,                 `f�)@ȵHPS!�?             :@       ������������������������       �                     0@        -       .                 �|�=@�z�G��?             $@        ������������������������       �                     �?        /       4                   @D@�<ݚ�?             "@       0       3                   �A@؇���X�?             @        1       2                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        5       6                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        9       V                    �?�)
;&��?>             W@        :       U                     �?�e����?            �C@       ;       T                   �H@��J�fj�?            �B@       <       Q                   @C@�g�y��?             ?@       =       >                   �4@�û��|�?             7@        ������������������������       �                     @        ?       P                 �̾w@�G�z��?             4@       @       M                    �?ҳ�wY;�?             1@       A       D                 �|�;@�q�q�?
             (@        B       C                 Ȉ�P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        E       L                   �A@�<ݚ�?             "@       F       K                 ��2>@�q�q�?             @        G       H                 `f&;@�q�q�?             @        ������������������������       �                     �?        I       J                 ���<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        N       O                   �7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        R       S                 ���X@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        W       f                  i?@�c�����?"            �J@        X       e                   @>@p�ݯ��?             3@       Y       d                   �J@�t����?
             1@       Z       c                 `f�;@X�<ݚ�?             "@       [       ^                 �|�?@����X�?             @        \       ]                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                   �C@z�G�z�?             @        ������������������������       �                     @        a       b                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        g       x                     �?@�0�!��?             A@       h       i                   �A@�n`���?             ?@        ������������������������       �                     "@        j       w                    �?���!pc�?             6@       k       v                    �?����X�?             5@       l       m                   �B@�z�G��?             4@        ������������������������       �                     @        n       u                 `f�K@@�0�!��?             1@       o       p                   �C@��S�ۿ?             .@       ������������������������       �                     "@        q       r                    �?r�q��?             @        ������������������������       �                     @        s       t                  x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        {       �                   �@@\�Yf�?�            �v@       |       �                    �?�8a�ME�?�            �s@        }       �                    �?@��Pl3�?<            @X@        ~       �                    �?     ��?             @@              �                    �?�>4և��?             <@       �       �                    �?�IєX�?             1@        ������������������������       �                      @        �       �                 �|�6@��S�ۿ?
             .@        ������������������������       �                     @        �       �                 ���@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?���|���?             &@        �       �                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?&����?(            @P@       �       �                 03�-@>���Rp�?%             M@       �       �                    �?�LQ�1	�?             G@       �       �                    �?8�Z$���?             :@       �       �                 ���@r�q��?             8@        ������������������������       �                     "@        �       �                   @@������?             .@       �       �                   �5@�q�q�?             "@        ������������������������       �                     �?        �       �                 �|=@      �?              @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        �       �                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y;@ףp=
�?             4@        ������������������������       �                     �?        �       �                  s�@�KM�]�?             3@        ������������������������       �                     @        �       �                    �?؇���X�?
             ,@       ������������������������       �8�Z$���?	             *@        ������������������������       �                     �?        �       �                 ��.@�q�q�?             (@        ������������������������       �                     @        �       �                 ��$1@և���X�?             @        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�nYU}�?�             k@       �       �                    @�C�F��?o            �e@       �       �                 �|�=@�R����?n            �e@       �       �                    �?*~k���?b            �b@        �       �                  s@�eP*L��?             6@        ������������������������       �                     @        �       �                    4@�q�q�?             2@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�;@d}h���?
             ,@       �       �                 pff@ףp=
�?             $@        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?x�]AgȽ?T             `@       �       �                    �?`Jj��?R             _@       �       �                 ���@�IєX�?N            �]@        �       �                   �5@����X�?             @        ������������������������       �                     @        �       �                 �&b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �0@���>4ֵ?I             \@        �       �                 pFD!@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        �       �                 @3�!@ 7���B�?E             [@       �       �                 @3�@������?6            �T@       �       �                 �?$@���J��?!            �I@        �       �                 ��@���N8�?             5@       ������������������������       �        	             1@        �       �                 �|Y8@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     >@        �       �                 pf� @��a�n`�?             ?@       �       �                   �4@�8��8��?             8@        �       �                   �2@����X�?             @        ������������������������       �                      @        �       �                 0S5 @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     1@        �       �                    8@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        �       �                 �Y�@z�G�z�?             @        ������������������������       �                      @        �       �                 pF�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@@8�A�0��?             6@       �       �                    �?      �?
             2@       �       �                    �?     ��?	             0@        ������������������������       �                     @        �       �                   �?@��
ц��?             *@        ������������������������       �                     @        �       �                 d�6@@���Q��?             $@       �       �                 ��I @և���X�?             @       �       �                 P�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �̜2@d}h���?             E@        �       �                    <@�	j*D�?             *@       �       �                 P�@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     H@        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  `l����??'��d�?G}g����?]AL� &�?|���?|���?�������?�������?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?��\V��?��FS���?�vV;��?���Tb*�?���̞?��g	�?AA�?~��}���?{�G�z�?\���(\�?�?�?              �?�������?�������?      �?      �?              �?      �?                      �?              �?�؉�؉�?ى�؉��?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?��]�`��?�T�6|��?���^B{�?/�����?��+��+�?�A�A�?      �?      �?      �?                      �?�������?�������?      �?              �?      �?��N��N�?�؉�؉�?      �?        ffffff�?333333�?              �?9��8���?�q�q�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?        ���7���?C���,�?�-��-��?�A�A�?�"�u�)�?к����?��{���?�B!��?8��Moz�?��,d!�?      �?        �������?�������?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        333333�?�������?              �?      �?                      �?      �?      �?              �?      �?              �?              �?        �V�9�&�?:�&oe�?^Cy�5�?Cy�5��?�������?�������?�q�q�?r�q��?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?              �?                      �?ZZZZZZ�?�������?�9�s��?�c�1��?      �?        F]t�E�?t�E]t�?�m۶m��?�$I�$I�?ffffff�?333333�?              �?ZZZZZZ�?�������?�������?�?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?              �?              �?              �?        p��.�^�?A�ME��?,��O[�?�O[h���?��4l7��?�n�'�i�?      �?      �?�m۶m��?�$I�$I�?�?�?              �?�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?]t�E]�?�������?�������?              �?      �?                      �?      �?        �����?�����?�i��F�?GX�i���?��Moz��?Y�B��?;�;��?;�;��?�������?UUUUUU�?      �?        wwwwww�?�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �������?UUUUUU�?              �?      �?              �?        �������?�������?      �?        �k(���?(�����?      �?        ۶m۶m�?�$I�$I�?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?        ӕ��te�?��Y�,j�?�L�w��?ȹ�. 6�?� �z�?��}���?��^x/�?�z=��?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        I�$I�$�?۶m۶m�?�������?�������?      �?      �?              �?      �?              �?              �?      �?      �?                      �?�?���?����?���{��?�B!��?�?�?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?%I�$I��?�m۶mۦ?      �?      �?      �?      �?      �?        	�%����?h/�����?p>�cp�?������?______�?�?��y��y�?�a�a�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �s�9��?�c�1Ƹ?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        颋.���?/�袋.�?      �?      �?      �?      �?              �?�;�;�?�؉�؉�?      �?        �������?333333�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?                      �?I�$I�$�?۶m۶m�?;�;��?vb'vb'�?F]t�E�?/�袋.�?      �?                      �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�F         D                    �?���Yb�?�           8�@               )                    �?&ջ�{��?]            @b@                                  �?JJ����?;            �W@                                   �?��hJ,�?             A@       ������������������������       �                     ;@                                �ܙH@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        	       
                   �2@      �?'             N@        ������������������������       �                     @                                     @����>4�?$             L@                                  @B@�ՙ/�?             5@                               ���<@      �?             0@        ������������������������       �                     @                                   �?�n_Y�K�?	             *@                               03SA@���Q��?             $@        ������������������������       �                     @                                @�6M@և���X�?             @        ������������������������       �                     @                                X�,@@      �?             @                               �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                �nc@�q�q�?             @        ������������������������       �                     �?                                �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               "                 �|Y=@�#-���?            �A@                !                   @@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        #       $                 ���@`2U0*��?             9@        ������������������������       �                     &@        %       (                 �|�=@@4և���?
             ,@       &       '                   @@      �?              @       ������������������������       �r�q��?             @        ������������������������       �                      @        ������������������������       �                     @        *       3                     @R�}e�.�?"             J@       +       ,                    �?z�G�z�?             >@       ������������������������       �                     4@        -       2                    �?���Q��?             $@       .       1                     �?�q�q�?             @       /       0                 �U�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        4       =                    �?���|���?
             6@        5       <                    �?և���X�?             ,@       6       9                    �?�eP*L��?             &@        7       8                   �-@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        :       ;                 �|Y3@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        >       C                 03�-@      �?              @       ?       B                    �?�q�q�?             @       @       A                 �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        E                       `f�S@��f
a�?r           ��@       F       �                 `f�$@�K�7���?]           Ȁ@        G       \                    �?��1��?�            �n@        H       S                   �6@�g�y��?             ?@        I       R                    �?r�q��?
             (@       J       O                    �?�<ݚ�?             "@       K       L                    �?؇���X�?             @        ������������������������       �                      @        M       N                   �3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       Q                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       Y                 ��@�d�����?             3@        U       V                 ���@�q�q�?             @        ������������������������       �                     �?        W       X                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       [                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ]       b                   �0@d��]a��?�            �j@        ^       _                 pf�@���!pc�?             &@        ������������������������       �                     @        `       a                 pFD!@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        c       l                    �?����p�?�            �i@        d       e                 ���@�>4և��?             <@        ������������������������       �                      @        f       g                 �|Y=@      �?
             4@        ������������������������       �                     @        h       k                 X��A@�t����?	             1@       i       j                    �?؇���X�?             ,@       ������������������������       �8�Z$���?             *@        ������������������������       �                     �?        ������������������������       �                     @        m       �                 �|�=@����!p�?u             f@       n       {                 �?$@ ,V�ނ�?V            �_@        o       x                 ���@�L���?            �B@       p       q                     @�g�y��?             ?@        ������������������������       �                     "@        r       s                  Md@���7�?             6@        ������������������������       �                     &@        t       u                    7@�C��2(�?             &@        ������������������������       �                     @        v       w                   �8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                 �|�;@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        |       �                    �?�x�E~�?;            @V@       }       �                    �?`���i��?:             V@       ~                        @3�@�D�e���?8            @U@        ������������������������       �                    �C@        �       �                   �;@�nkK�?             G@       �       �                   �9@�>����?             ;@       �       �                   �3@ ��WV�?             :@        �       �                   �2@�C��2(�?             &@        ������������������������       �                     @        �       �                 0S5 @؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @@@ףp=
�?             I@        �       �                 �?�@�	j*D�?             *@        ������������������������       �                     @        �       �                    ?@X�<ݚ�?             "@        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��I @և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                      @�?�|�?            �B@        ������������������������       �                     @        �       �                   �C@г�wY;�?             A@       �       �                   @C@�IєX�?             1@       ������������������������       �        
             .@        ������������������������       �      �?              @        ������������������������       �        	             1@        �       �                    �?��c���?�            0r@        �       �                    �?ڷv���?I            �\@        �       �                    �?Hm_!'1�?            �H@        ������������������������       �                     �?        �       �                    �?      �?             H@       �       �                     @ �Cc}�?             <@       �       �                     �?$�q-�?             :@        ������������������������       �                     @        �       �                   �A@�C��2(�?             6@       �       �                   �9@�IєX�?
             1@        �       �                   �'@؇���X�?             @        ������������������������       �                     @        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                     @8�A�0��?*            �P@        �       �                     �?�}�+r��?             3@        ������������������������       �                     @        �       �                    �?��S�ۿ?             .@        �       �                    B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    �?��k=.��?            �G@        ������������������������       �                      @        �       �                   @1@���V��?            �F@        �       �                    �?���|���?             &@       �       �                    D@����X�?             @       �       �                 �|�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @l��\��?             A@        �       �                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @ 7���B�?             ;@       ������������������������       �                     7@        �       �                   @D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?��|���?t             f@       �       �                    �?H%u��?T            @_@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 `fF:@�S#א��?N            @]@       �       �                    4@����p�?+             Q@        �       �                    &@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                     @����˵�?$            �M@       �       �                   �*@���.�6�?             G@       �       �                 `f�)@ܷ��?��?             =@        ������������������������       �                     @        �       �                   �A@�LQ�1	�?             7@       �       �                    @@d}h���?             ,@       ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     "@        ������������������������       �                     1@        ������������������������       �                     *@        �                         �Q@Jm_!'1�?#            �H@       �                          �?r�q��?"             H@       �                             @t/*�?!            �G@       �       �                   �;@"pc�
�?             F@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@�p ��?            �D@        �       �                    K@     ��?             0@       �       �                   `G@�eP*L��?             &@       �       �                   @>@      �?              @       �       �                 `f�;@؇���X�?             @       �       �                 �|�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@`2U0*��?             9@       ������������������������       �                     1@        �       �                 `�iJ@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��[�8��?             �I@                                +@J�8���?             =@        ������������������������       �                     $@        ������������������������       �                     3@                                 @���7�?             6@       	      
                   �?      �?
             0@       ������������������������       �                     *@                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�>4և��?             <@                                M@H%u��?             9@                              �k@�8��8��?             8@                               @E@�nkK�?             7@       ������������������������       �                     3@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  �\	��`�?�F�+J>�?����?�?~���?��
br�?x6�;��?�������?KKKKKK�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?      �?              �?n۶m۶�?I�$I�$�?�<��<��?�a�a�?      �?      �?      �?        ى�؉��?;�;��?�������?333333�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �A�A�?_�_�?�������?�������?      �?                      �?���Q��?{�G�z�?      �?        n۶m۶�?�$I�$I�?      �?      �?�������?UUUUUU�?      �?              �?        �;�;�?'vb'vb�?�������?�������?              �?333333�?�������?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?              �?        F]t�E�?]t�E]�?۶m۶m�?�$I�$I�?t�E]t�?]t�E�?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?.rt�"G�?�9�q�?N��B�1�?�	��9�?�+Q���?,Q��+�?�B!��?��{���?UUUUUU�?�������?�q�q�?9��8���?�$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?      �?      �?              �?      �?                      �?Cy�5��?y�5���?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        �؉�؉�?;�;��?              �?      �?        �"�{(R�?��V!�n�?F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?        �������?�����Ҳ?�$I�$I�?�m۶m��?      �?              �?      �?              �?<<<<<<�?�?۶m۶m�?�$I�$I�?;�;��?;�;��?      �?              �?        /�袋.�?]t�E�?�뺮��?EQEQ�?}���g�?L�Ϻ��?��{���?�B!��?      �?        �.�袋�?F]t�E�?      �?        ]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?����G�?p�\��?F]t�E�?F]t�E�???????�?�?      �?        �Mozӛ�?d!Y�B�?�Kh/��?h/�����?O��N���?;�;��?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?                      �?      �?              �?              �?        �������?�������?vb'vb'�?;�;��?      �?        r�q��?�q�q�?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?�������?333333�?      �?        *�Y7�"�?к����?      �?        �?�?�?�?      �?              �?      �?      �?        �&�.9�?��ǿ���?]R�0��?A�V���?9/���?Y�Cc�?      �?              �?      �?۶m۶m�?%I�$I��?;�;��?�؉�؉�?              �?F]t�E�?]t�E�?�?�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?      �?      �?      �?                      �?              �?颋.���?/�袋.�?(�����?�5��P�?              �?�?�������?      �?      �?              �?      �?                      �?g���Q��?br1���?              �?[�[��?�>�>��?]t�E]�?F]t�E�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        ------�?�������?�m۶m��?�$I�$I�?      �?                      �?	�%����?h/�����?      �?              �?      �?              �?      �?        F]t�E�?颋.���?)\���(�?���Q��?      �?      �?      �?                      �?��+��+�?�꡾?�������?�����Ҳ?9��8���?�q�q�?              �?      �?        W'u_�?��/���?���7���?Y�B��?��=���?a���{�?      �?        ��Moz��?Y�B��?I�$I�$�?۶m۶m�?      �?              �?      �?      �?              �?              �?        ����X�?������?�������?UUUUUU�?�;����?W�+���?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?Q��+Q�?��+Q��?      �?      �?t�E]t�?]t�E�?      �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?                      �?              �?      �?        ���Q��?{�G�z�?      �?              �?      �?              �?      �?              �?              �?                      �?�?�������?�rO#,��?|a���?              �?      �?        �.�袋�?F]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?���Q��?)\���(�?UUUUUU�?UUUUUU�?d!Y�B�?�Mozӛ�?              �?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bub�0>     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM	hvh)h,K ��h.��R�(KM	��h}�B@B         l                 ��%@�*���?�           8�@                                   /@,PY��?�             v@        ������������������������       �                     @                                ���@j�q����?�            �u@        ������������������������       �                    �E@               3                 P�*@�A��t��?�            0s@               2                 �|Y>@J��D��?A             [@              1                    �?���Q �?8            �X@       	       
                 ��@r�qG�?7             X@        ������������������������       �                     �?                                   �?�|R���?6            �W@                                  �3@���B���?             :@                                �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�LQ�1	�?             7@                                  8@�C��2(�?             6@        ������������������������       �                     "@                                ��@8�Z$���?	             *@                               ���@�C��2(�?             &@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               $                   �<@�㙢�c�?&            @Q@               #                   �6@�C��2(�?            �@@                                  �3@�S����?
             3@        ������������������������       �                      @        !       "                    �?���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        %       .                    �?      �?             B@       &       '                 ���@z�G�z�?             9@        ������������������������       �                      @        (       )                 �|Y=@�t����?             1@        ������������������������       �                     �?        *       +                 ���@      �?
             0@        ������������������������       ����Q��?             @        ,       -                 �Y�@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �      �?              @        /       0                 ��,@���|���?             &@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �        	             $@        4       i                    �?ȭ^���?x            �h@       5       <                 �?�@��ɉ�?v            `h@        6       ;                 �̌@�L#���?)            �P@        7       8                 �|Y=@���y4F�?             3@       ������������������������       �        
             *@        9       :                 ��]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     H@        =       B                     @     ��?M             `@        >       A                   �J@�+e�X�?             9@       ?       @                    �?�����?             3@        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @        C       N                 @3�@�v�G���??            �Y@        D       G                    �?      �?             0@        E       F                   �9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        H       I                    :@���|���?             &@        ������������������������       �                     @        J       K                   �?@և���X�?             @        ������������������������       �                     �?        L       M                   �A@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        O       V                   �:@�=C|F�?4            �U@        P       U                   �3@`Ӹ����?            �F@        Q       T                 0S5 @�����?
             5@        R       S                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     8@        W       X                   �;@d}h���?             E@        ������������������������       �                     @        Y       h                   �?@8�Z$���?            �C@       Z       [                 ��) @      �?             8@       ������������������������       �        	             &@        \       ]                   �<@��
ц��?             *@        ������������������������       �                     @        ^       c                 P�*"@���Q��?             $@        _       `                 pf� @z�G�z�?             @        ������������������������       �                      @        a       b                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       e                 ���"@���Q��?             @        ������������������������       �                      @        f       g                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             .@        j       k                   �#@      �?             @        ������������������������       �                      @        ������������������������       �                      @        m       �                  x#J@��d���?�            Pv@       n       �                    �?~���n��?�            Pp@        o       �                    @t�I��n�?R            @]@       p       u                    @f�����?N            �[@        q       r                    @�}�+r��?             3@       ������������������������       �        
             0@        s       t                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       �                     @ �&�T�?B             W@       w       �                   �H@�j��b�?(            �M@       x       �                    �?,�+�C�?%            �K@       y       z                     �?<���D�?            �@@        ������������������������       �                     @        {       �                   �7@8�Z$���?             :@       |       �                    �?������?             .@       }       �                    :@d}h���?             ,@        ~                           �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ףp=
�?	             $@        ������������������������       �                     �?        �       �                   �*@�����H�?             "@       �       �                 `f�)@؇���X�?             @        ������������������������       �                     �?        �       �                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     6@        �       �                 03�9@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?4���C�?            �@@       �       �                 ��.@\X��t�?             7@       �       �                    �?�	j*D�?
             *@        �       �                 �|Y6@և���X�?             @       �       �                   �,@      �?             @        ������������������������       �                      @        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �*@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 �|Y>@r�q��?             @        ������������������������       �                     @        �       �                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���0@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    @�q�q�?g             b@       �       �                    !@�θ�?^            @`@        ������������������������       �                     $@        �       �                 �&@r�q��?W             ^@        ������������������������       �                     �?        �       �                     �?�?��,�?V            �]@        �       �                 ��";@���j��?             G@        �       �                 ��$:@և���X�?
             ,@        ������������������������       �                     @        �       �                   �J@���!pc�?             &@       �       �                   @G@�����H�?             "@       �       �                    D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?     ��?             @@       �       �                 ���=@�����?             5@        ������������������������       �                     $@        �       �                 p�i@@"pc�
�?             &@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@���!pc�?	             &@        ������������������������       �                      @        �       �                 �|Y>@�����H�?             "@        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �*@�F��O�?8            @R@        �       �                   �@@�㙢�c�?             7@       ������������������������       �        
             (@        �       �                   �)@���|���?	             &@        ������������������������       �                      @        �       �                   �A@X�<ݚ�?             "@        ������������������������       �      �?             @        �       �                   @D@z�G�z�?             @        ������������������������       �                      @        �       �                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`2U0*��?%             I@       �       �                 ��.@`Ql�R�?"            �G@        �       �                     @$�q-�?
             *@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        �                          @     ��?B             X@       �       �                    �?�n`���??            @W@       �       �                   �5@f>�cQ�?-            �N@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?$�q-�?'             J@       �       �                      @�IєX�?&            �I@       �       �                   �B@ �q�q�?#             H@       �       �                    �?�IєX�?             A@       ������������������������       �                     <@        �       �                    �?�q�q�?             @       �       �                 X�,@@      �?             @       �       �                 p"�b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 �7@     ��?             @@                                 �?�C��2(�?             &@                                �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�ՙ/�?             5@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM	KK��h^�B�  P�D��n�?auv�4"�?�s�f���?-1>e�9�?              �?=
ףp=�?
ףp=
�?      �?        �M��n�?M�ɺ`D�?�^B{	��?_B{	�%�?9/����?����>4�?�������?�������?              �?&N��[��?�c�H;�?ى�؉��?��؉���?UUUUUU�?UUUUUU�?              �?      �?        Y�B��?��Moz��?F]t�E�?]t�E�?              �?;�;��?;�;��?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?        �7��Mo�?d!Y�B�?]t�E�?F]t�E�?(������?^Cy�5�?      �?        F]t�E�?t�E]t�?              �?      �?              �?              �?      �?�������?�������?      �?        �������?�������?              �?      �?      �?�������?333333�?]t�E�?F]t�E�?      �?              �?      �?]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?              �?        �|i�0V�?�Zv<��?�����?�����?��@���?g��1��?6��P^C�?(������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?             @�?      �?R���Q�?���Q��?Q^Cy��?^Cy�5�?              �?      �?              �?        C���?��O �?      �?      �?333333�?�������?      �?                      �?]t�E]�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?      �?�C��:��?J��/�??�>��?l�l��?=��<���?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        I�$I�$�?۶m۶m�?              �?;�;��?;�;��?      �?      �?      �?        �;�;�?�؉�؉�?      �?        �������?333333�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        ^9�]9��?Q�Q��?M�s���?e�� 3�?���?�s?�s?�?���+c��?�5'��?(�����?�5��P�?              �?UUUUUU�?UUUUUU�?      �?                      �?���,d�?��7��M�?��/���?�N��?��)A��?�}��7��?|���?|���?              �?;�;��?;�;��?�?wwwwww�?۶m۶m�?I�$I�$�?      �?      �?              �?      �?        �������?�������?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?      �?                      �?      �?                      �?              �?      �?      �?              �?      �?        m��&�l�?'�l��&�?��Moz��?!Y�B�?vb'vb'�?;�;��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?              �?      �?        �������?�������?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?�������?�������?              �?      �?              �?        UUUUUU�?�������?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?              �?����?��o��o�?ozӛ���?!Y�B�?۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?�q�q�?�q�q�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?=��<���?�a�a�?      �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �իW�^�?�P�B�
�?�7��Mo�?d!Y�B�?      �?        ]t�E]�?F]t�E�?      �?        r�q��?�q�q�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���Q��?{�G�z�?}g���Q�?W�+�ɕ?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?�c�1��?�9�s��?�u�y���?��!XG�?r�q��?�q�q�?              �?      �?        ;�;��?�؉�؉�?�?�?UUUUUU�?�������?�?�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?F]t�E�?]t�E�?�������?�������?      �?                      �?              �?�a�a�?�<��<��?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM	hvh)h,K ��h.��R�(KM	��h}�B@B         p                     @���%&�?�           8�@               '                 �|Y=@N�ec�?�            ps@               
                 ��*@"��$�?G            �[@               	                    �?      �?             8@                                   �?"pc�
�?             &@                               `f�)@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@               "                 `fmj@�N��D�?6            �U@                                  �?���(\��?2             T@                                  6@�C��2(�?)            �P@                                   9@���|���?             &@       ������������������������       �                     @                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?h㱪��?#            �K@       ������������������������       �                    �B@                                    �?�����H�?
             2@                                  5@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?d}h���?	             ,@                                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                !                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        #       &                 0U�o@և���X�?             @       $       %                    5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        (       9                    �?4��@���?�             i@        )       ,                    �?�nkK�?1            @Q@        *       +                 03�=@`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        -       6                    L@���7�?             F@       .       /                   �B@��Y��]�?            �D@       ������������������������       �                     8@        0       5                    -@�IєX�?             1@        1       2                   �'@�q�q�?             @        ������������������������       �                     �?        3       4                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        7       8                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        :       o                   �J@��ׂ�?Z            ``@       ;       n                 p�w@������?F            @Z@       <       a                   �G@��z6��?D             Y@       =       >                   �)@� ���?6            @S@        ������������������������       �        	             ,@        ?       `                   �F@��s����?-            �O@       @       [                    �?�T`�[k�?(            �J@       A       L                    �?��Q���?             D@        B       K                    �?     ��?
             0@       C       J                    C@�q�q�?	             .@       D       I                 ��2>@����X�?             ,@        E       H                 ���<@      �?              @       F       G                 ��";@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        M       Z                    �?      �?             8@       N       W                   @D@���!pc�?             6@       O       V                 `f�<@@�0�!��?             1@       P       U                 `fF:@���!pc�?             &@       Q       T                 `fv3@z�G�z�?             $@       R       S                 �|�=@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                     �?���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                      @        \       ]                   �B@$�q-�?             *@        ������������������������       �                     @        ^       _                 03�U@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        b       c                 `f4@
;&����?             7@        ������������������������       �                     @        d       i                    �?     ��?	             0@        e       f                    �?�q�q�?             @        ������������������������       �                      @        g       h                 ���X@      �?             @       ������������������������       �                      @        ������������������������       �                      @        j       k                 ���E@ףp=
�?             $@       ������������������������       �                      @        l       m                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        q                          @z6�>��?            y@       r       s                 ���@�o6�
�?�            �x@        ������������������������       �                     ;@        t                          @.�6�G,�?�             w@       u       �                    �?H?�߽��?�            �v@        v       �                    �?�\��N��?H            �\@        w       |                    �?,���i�?            �D@       x       {                 ���@      �?             @@        y       z                 0��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        }       ~                    @X�<ݚ�?             "@        ������������������������       �                      @               �                  S�2@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                 ���&@�q�q�?             @        ������������������������       �                     �?        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @:PZ(8?�?-            @R@        �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ,@�t����?)             Q@        ������������������������       �                     $@        �       �                   �"@J�8���?$             M@        �       �                    @�ՙ/�?             5@       �       �                    ;@���Q��?             4@       �       �                    �?������?
             .@       �       �                 pf� @d}h���?	             ,@       �       �                   �7@�C��2(�?             &@        ������������������������       �                     @        �       �                 �&B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?� @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�1@��G���?            �B@       �       �                    �?�X����?             6@       �       �                     @ҳ�wY;�?             1@       �       �                   �3@������?
             .@        ������������������������       �                     �?        �       �                   �0@d}h���?	             ,@       �       �                 �|�;@8�Z$���?             *@        ������������������������       �                      @        �       �                 ���.@���Q��?             @       �       �                    �?      �?             @       �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                 ��@H%u��?�            @o@        ������������������������       �                     @        �       �                    #@0�v����?�            �n@        �       �                     @     ��?             0@        ������������������������       �                     @        �       �                    @ףp=
�?             $@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 ���A@      �?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?,���>�?�            �l@        �       �                 03�-@д>��C�?'             M@       �       �                 �|Y=@ףp=
�?              I@        �       �                   �<@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y?@��p\�?            �D@       �       �                    �?ܷ��?��?             =@       �       �                 ���@�����H�?             ;@        ������������������������       �                     @        �       �                 P�J@؇���X�?             5@       �       �                 ���@R���Q�?             4@        �       �                    �?�����H�?             "@       ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �"pc�
�?             &@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                 ��.@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �                         @@@���y�?p            �e@       �                          �?D��*�4�?\            @a@       �                          �?�[|x��?U            �_@       �       �                 �!&B@�H�@=��?M            �[@       �       �                 �|�=@ �h�7W�?J            �Z@       �       �                 @3�@��8�$>�?C            @X@       ������������������������       �        $             H@        �       �                 @�!@Hm_!'1�?            �H@       �       �                   � @PN��T'�?             ;@       �       �                 0S5 @�r����?             .@       �       �                   �3@؇���X�?             ,@        �       �                    1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �7@r�q��?             (@       ������������������������       �                      @        �       �                 �|Y<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        �       �                   �?@�<ݚ�?             "@       �       �                   �>@���Q��?             @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ;@z�G�z�?             @        ������������������������       �                      @                                  >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     (@        ������������������������       �                    �A@                               �:@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM	KK��h^�B�  �g *��?�0���M�?�p�X��?�G�S6�?Nq��$�?�~G����?      �?      �?F]t�E�?/�袋.�?�q�q�?9��8���?              �?      �?                      �?      �?        �2)^ �?�~�u�7�?�����̼?ffffff�?F]t�E�?]t�E�?F]t�E�?]t�E]�?              �?�������?�������?              �?      �?        ��)A��?־a���?              �?�q�q�?�q�q�?�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?I�$I�$�?�q�q�?�q�q�?      �?                      �?�������?333333�?              �?      �?        �$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?�(\����?�G�z�?d!Y�B�?�Mozӛ�?{�G�z�?���Q��?      �?                      �?F]t�E�?�.�袋�?������?8��18�?              �?�?�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?w�_�	)�?#����[�?wwwwww�?�?�p=
ף�?q=
ףp�?L�S�?��O����?      �?        z��y���?�a�a�?���!5��?"5�x+��?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?      �?�������?�������?              �?      �?                      �?      �?                      �?      �?              �?      �?F]t�E�?t�E]t�?ZZZZZZ�?�������?F]t�E�?t�E]t�?�������?�������?�m۶m��?�$I�$I�?              �?      �?              �?                      �?      �?        �������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?        �؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?                      �?      �?        Y�B��?�Mozӛ�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?              �?      �?        ���(\��?��(\���?�}z)@w�?	Z�"�?      �?        ���7���?C���,�?h�h��?`��_���?�5��P�?y�5���?8��18�?�����?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�W�^�z�?�P�B�
�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        �rO#,��?|a���?�a�a�?�<��<��?�������?333333�?�?wwwwww�?۶m۶m�?I�$I�$�?F]t�E�?]t�E�?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?      �?                      �?              �?#�u�)��?v�)�Y7�?�E]t��?]t�E]�?�������?�������?wwwwww�?�?              �?I�$I�$�?۶m۶m�?;�;��?;�;��?      �?        333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?              �?              �?�������?�������?              �?      �?              �?        )\���(�?���Q��?              �?������?��1����?      �?      �?              �?�������?�������?�������?�������?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        ���e�:�?s�X�*�?a���{�?|a���?�������?�������?9��8���?�q�q�?      �?                      �?�]�ڕ��?��+Q��?��=���?a���{�?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?333333�?333333�?�q�q�?�q�q�?�������?UUUUUU�?      �?        /�袋.�?F]t�E�?      �?              �?              �?              �?      �?              �?333333�?�������?              �?      �?      �?      �?                      �?�mNWy&�?�'�j��?ہ�v`��?)�3J���?]�u]�u�?EQEQ�?��+c��?q��$�?��sHM0�?"5�x+��?�Q�/��?����?      �?        Y�Cc�?9/���?&���^B�?h/�����?�������?�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?UUUUUU�?      �?              �?      �?              �?      �?              �?        9��8���?�q�q�?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�C         \                    �?�s�ˈ.�?�           8�@               U                 p�H@�d�����?�            �l@              4                    �?Ҙ$�Ų�?k            �d@                                   @�<ݚ�?=            �X@               
                    �?�(\����?             D@                                 �J@�nkK�?             7@       ������������������������       �                     4@               	                 `f�2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@                                   �?:���W�?#            �M@                                   �?�+e�X�?             9@                                H�%@���Q��?             $@        ������������������������       �                     @                                03�-@z�G�z�?             @        ������������������������       �                     @                                �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                X�,A@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @               /                    �?�ʻ����?             A@              .                    �?*;L]n�?             >@                                  '@П[;U��?             =@        ������������������������       �                     @                                  �4@      �?             :@        ������������������������       �                     @               )                 `��!@\X��t�?             7@              (                    C@������?	             .@               !                 P�@d}h���?             ,@        ������������������������       �                     @        "       '                 �|Y>@      �?              @       #       &                 �|�;@      �?             @       $       %                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        *       +                    ;@      �?              @       ������������������������       �                     @        ,       -                   �@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                    @      �?             @        ������������������������       �                     �?        2       3                 ��l4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        5       <                     @�'�=z��?.            �P@        6       9                    6@؇���X�?             5@        7       8                 ��m1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        :       ;                   �B@�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        =       @                    �?f.i��n�?            �F@        >       ?                 ��.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        A       J                 03�1@��Sݭg�?            �C@        B       I                    �?�q�q�?             (@       C       H                 ��Y.@���Q��?             $@       D       G                    �?z�G�z�?             @       E       F                    6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        K       P                    @�>����?             ;@       L       O                 ���4@���7�?             6@        M       N                 03C3@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             3@        Q       R                 ��T?@z�G�z�?             @        ������������������������       �                      @        S       T                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        V       [                 ���Q@$Q�q�?+            �O@        W       X                    �?�J�4�?             9@       ������������������������       �                     3@        Y       Z                 ���P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     C@        ]       �                    �?���A�
�?*           0~@        ^       k                 ��K.@N��c��?1            @S@        _       d                   �6@������?            �D@        `       a                    �?      �?             @        ������������������������       �                     �?        b       c                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                 �|=@�?�|�?            �B@        ������������������������       �                     &@        g       j                   @@ ��WV�?             :@       h       i                 ���@�C��2(�?             &@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     .@        l       w                    �?b�2�tk�?             B@       m       r                 �|Y<@�z�G��?             4@        n       q                    9@����X�?             @        o       p                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        s       v                   �F@$�q-�?
             *@        t       u                 X�,@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        x                           �?      �?             0@       y       |                 ��G@և���X�?
             ,@        z       {                 ��3@      �?              @        ������������������������       �                     @        ������������������������       �                     @        }       ~                 ���X@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �/@|g�&��?�            `y@       �       �                    �?<N_�U��?�            �p@       �       �                 �?�@     �?�             p@        �       �                     @������?M            �^@        ������������������������       �                     &@        �       �                    �?�h����?E             \@        �       �                  ��@8�Z$���?             *@        ������������������������       �                      @        �       �                    �?"pc�
�?	             &@       �       �                 �|Y=@�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��(@      �?              @       ������������������������       �r�q��?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �7@��:x�ٳ?:            �X@        ������������������������       �                     A@        �       �                 �Yu@����?&            @P@       �       �                 �&B@(N:!���?            �A@       �       �                   �8@`Jj��?             ?@        �       �                 �&b@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     >@        �       �                   �0@���H��?N            �`@        �       �                 �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �*@ ����?L            @`@       �       �                   �A@���5��?D            �\@       �       �                   �<@8�Z$���?7            �V@       �       �                   �3@$�q-�?             J@        �       �                     @������?	             .@        �       �                    &@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        �       �                   �1@���!pc�?             &@        ������������������������       �                     @        �       �                 0S5 @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �B@        �       �                 ��)"@��Sݭg�?            �C@       �       �                   �?@�KM�]�?             3@       �       �                   �>@8�Z$���?             *@       �       �                 �|Y=@�8��8��?
             (@        ������������������������       �                     �?        �       �                 ��) @�C��2(�?	             &@       ������������������������       �                     "@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@���Q��?             4@        ������������������������       �                     @        �       �                   �@@�t����?             1@       �       �                    $@�θ�?	             *@        �       �                   �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �      �?             @        ������������������������       �                     7@        ������������������������       �                     0@        �       �                    �?���|���?             &@       �       �                     @X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �*@      �?              @        �       �                 xFT$@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @4kMU*m�?X            `a@        �       �                   �;@������?             .@        ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        �                          �?���b��?P             _@       �       �                    �? �&�T�?:             W@       �       �                     @���3�E�?$             J@       �       �                 ��$:@�*/�8V�?             �G@        ������������������������       �        	             .@        �       �                   �>@      �?             @@       �       �                 `fF<@�t����?             1@       �       �                    K@      �?             $@       �       �                 03k:@����X�?             @        ������������������������       �                     �?        �       �                 �|�<@�q�q�?             @        ������������������������       �                      @        �       �                 X��B@      �?             @        ������������������������       �                     �?        �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        �       �                 �|�>@���Q��?             @       �       �                 �T�C@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             D@       �       �                  x#J@r٣����?            �@@       ������������������������       �        
             1@        �       �                    F@      �?             0@       �       �                 `f�K@�q�q�?             (@       �       �                    7@      �?              @        ������������������������       �                     @        �       �                 `�iJ@z�G�z�?             @        ������������������������       �                      @        �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�:@����X�?             @        ������������������������       �                     @                                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 @      �?             @@                                �?`Jj��?             ?@                                 @�X�<ݺ?             2@        ������������������������       �                     @              
                   @@4և���?	             ,@             	                   0@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  ��0Ȍ��?��o��?y�5���?Cy�5��?��[���?$�:R�#�?�q�q�?9��8���?�������?333333�?d!Y�B�?�Mozӛ�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?A�Iݗ��?_[4��?���Q��?R���Q�?�������?333333�?              �?�������?�������?      �?              �?      �?              �?      �?        �?�������?              �?      �?        <<<<<<�?�������?�������?""""""�?��=���?�{a���?              �?      �?      �?      �?        ��Moz��?!Y�B�?�?wwwwww�?۶m۶m�?I�$I�$�?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        |��|�?|���?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        �?�?              �?      �?        �`�`�?�>�>��?UUUUUU�?UUUUUU�?      �?                      �?�|˷|��?�i�i�?UUUUUU�?UUUUUU�?�������?333333�?�������?�������?      �?      �?              �?      �?              �?                      �?              �?�Kh/��?h/�����?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        AA�?~��}���?{�G�z�?�z�G��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?��9��?7�5���?�����?5�wL��?�|����?������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        *�Y7�"�?к����?      �?        O��N���?;�;��?]t�E�?F]t�E�?      �?              �?      �?      �?        �8��8��?9��8���?ffffff�?333333�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?�؉�؉�?;�;��?�������?�������?      �?                      �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?              �?        ��v���?��%f-�?���F��?�!�c��?     @�?      �?p>�cp�?������?      �?        �$I�$I�?۶m۶m�?;�;��?;�;��?      �?        /�袋.�?F]t�E�?9��8���?�q�q�?              �?      �?      �?�������?UUUUUU�?      �?              �?        
�����?[�R�֯�?      �?        ~�~��? �����?|�W|�W�?�A�A�?���{��?�B!��?333333�?�������?      �?                      �?      �?              �?      �?              �?      �?              �?        h	&�?���̾?UUUUUU�?UUUUUU�?              �?      �?        �ȍ�ȍ�?�����?�}��?��Gp�?;�;��?;�;��?�؉�؉�?;�;��?wwwwww�?�?      �?      �?      �?      �?      �?        F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        �|˷|��?�i�i�?�k(���?(�����?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?                      �?      �?        333333�?�������?              �?�������?�������?ى�؉��?�؉�؉�?      �?      �?              �?      �?              �?              �?      �?      �?              �?        ]t�E]�?F]t�E�?r�q��?�q�q�?              �?      �?      �?�������?333333�?      �?                      �?      �?              �?        �R��u@�??ZMB�?�?wwwwww�?              �?      �?      �?              �?      �?        !�B�?�{����?��7��M�?���,d�?O��N���?b'vb'v�?�٨�l��?AL� &W�?      �?              �?      �?�������?�������?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?>���>�?|���?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?���{��?�B!��?��8��8�?�q�q�?      �?        n۶m۶�?�$I�$I�?�q�q�?�q�q�?              �?      �?              �?        �؉�؉�?;�;��?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK���h}�B@?         b                    �?��eC~�?�           8�@               ]                 p�H@������?�            `n@              D                    �?�H�]�r�?p            @e@              	                 ��@r�0p�?F            �Z@                                   �?P���Q�?             4@       ������������������������       �        	             ,@                                ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        
                            @��V#�?8            �U@                                   L@>A�F<�?             C@                                  �?     ��?             @@        ������������������������       �                     @                                `f�)@�����H�?             ;@        ������������������������       �                     &@                                   �?     ��?             0@                                  :@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@                                   <@      �?             @                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                `f�2@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @               7                 �|�<@     ��?              H@              ,                 Ь�!@�5��?             ;@              #                   �6@���Q��?             .@               "                 �&B@�<ݚ�?             "@                !                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        $       %                 �&B@�q�q�?             @        ������������������������       �                     �?        &       '                   �9@���Q��?             @        ������������������������       �                      @        (       )                   �@�q�q�?             @        ������������������������       �                     �?        *       +                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -       0                    �?r�q��?	             (@        .       /                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        1       6                 ��.@�����H�?             "@       2       3                   �-@z�G�z�?             @        ������������������������       �                      @        4       5                 �yG(@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        8       =                 �|Y>@���N8�?             5@       9       :                    �?@4և���?             ,@       ������������������������       �                     $@        ;       <                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        >       A                    @@և���X�?             @        ?       @                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        B       C                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        E       J                    �?      �?*             P@        F       I                    �?���Q��?	             .@       G       H                 `�@1@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        K       L                    @Rg��J��?!            �H@        ������������������������       �                     @        M       N                    (@��6���?             E@        ������������������������       �                      @        O       P                   �:@�ʻ����?             A@        ������������������������       �        
             &@        Q       \                     @�LQ�1	�?             7@       R       [                    @X�<ݚ�?
             2@       S       T                   �?@��.k���?	             1@        ������������������������       �                     @        U       V                     @�q�q�?             (@        ������������������������       �                     @        W       X                    �?      �?              @        ������������������������       �                      @        Y       Z                 ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                    !@��pBI�?0            @R@        ������������������������       �                     �?        `       a                    @�k~X��?/             R@       ������������������������       �        .            �Q@        ������������������������       �                     �?        c       n                    @K�(i�?"           @}@        d       i                    �?8����?             7@       e       f                     @�q�q�?             (@       ������������������������       �                     @        g       h                 �y�-@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        j       k                     @"pc�
�?             &@       ������������������������       �                     @        l       m                 pf�@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        o       �                    �?4�<����?           �{@        p       {                 P�J.@����X�?4             U@        q       r                   @@     ��?             @@       ������������������������       �                     1@        s       z                 �(@z�G�z�?             .@        t       y                 �y�#@և���X�?             @       u       x                 �� @z�G�z�?             @       v       w                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        |       �                    �?�E��
��?              J@       }       �                   �H@j���� �?            �I@       ~       �                     @      �?             E@              �                     �?��%��?            �B@       �       �                   �8@*;L]n�?             >@        �       �                  D�U@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             8@       �       �                 �ܵ<@      �?             4@        ������������������������       �                      @        �       �                    �?r�q��?
             2@       �       �                 `f�A@      �?             (@        ������������������������       �                     @        �       �                 @�6M@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 @��v@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                 `ff:@���5���?�            �v@       �       �                    �?��S�jC�?�            pr@       �       �                    )@(�s���?�            �o@        ������������������������       �                      @        �       �                   @E@ ��GS=�?�            @o@       �       �                   �D@�IєX�?�            �k@       �       �                 ���@�X�<ݺ?�             k@        ������������������������       �                    �C@        �       �                 �?$@ ,��-�?i             f@        �       �                   �;@�㙢�c�?             7@        ������������������������       �                     @        �       �                    �?������?
             1@       �       �                 �|Y=@d}h���?             ,@        ������������������������       �                      @        ������������������������       ��8��8��?             (@        �       �                 �|Y?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@�kb97�?[            @c@        ������������������������       �                    �A@        �       �                   �3@T(y2��?C            �]@        �       �                   �1@��2(&�?             6@        ������������������������       �                     @        �       �                 0S5 @z�G�z�?	             .@        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     &@        �       �                    �?h�a��?7            @X@       �       �                 �|�=@ rpa�?5            @W@       �       �                 @3�!@��v$���?!            �N@        �       �                 pf� @�nkK�?             7@       ������������������������       �        
             4@        �       �                    8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     C@        �       �                   �?@      �?             @@        �       �                     @�<ݚ�?             "@        ������������������������       �                     @        �       �                 @3�@      �?             @        ������������������������       �                     �?        �       �                 �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �@@���}<S�?             7@        ������������������������       �                     "@        �       �                     @؇���X�?	             ,@       �       �                   �3@؇���X�?             @       �       �                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 @3�@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���%@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     =@        �       �                     @ qP��B�?            �E@        ������������������������       �                      @        �       �                   �/@��?^�k�?            �A@       ������������������������       �                     2@        �       �                    )@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    �?:ɨ��?-            �P@       �       �                    �?���Q��?              I@       �       �                     �?��.k���?             A@       �       �                   �>@X�<ݚ�?             ;@       �       �                    R@����X�?             5@       �       �                   @=@�q�q�?             2@       �       �                 �|�<@���Q��?             $@        ������������������������       �                     �?        �       �                 `f�;@�q�q�?             "@       �       �                 �|�?@      �?              @        ������������������������       �                     @        �       �                   �J@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�>@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��9L@      �?
             0@       �       �                   �C@ףp=
�?             $@        ������������������������       �                     @        �       �                    G@�q�q�?             @       �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �D@      �?             @       �       �                     �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        �t�b��     h�h)h,K ��h.��R�(KK�KK��h^�B�  ���Kkz�?�fh)�?{	�%���?B{	�%��?�������?�������?oe�Cj��?HM0��>�?�������?ffffff�?              �?UUUUUU�?�������?              �?      �?        6eMYS��?eMYS֔�?Cy�5��?������?      �?      �?              �?�q�q�?�q�q�?              �?      �?      �?UUUUUU�?�������?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?h/�����?/�����?�������?333333�?�q�q�?9��8���?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��y��y�?�a�a�?�$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?333333�?�������?]t�E�?t�E]t�?      �?                      �?      �?        ��S�r
�??4և���?              �?b�a��?=��<���?      �?        <<<<<<�?�������?              �?Nozӛ��?d!Y�B�?r�q��?�q�q�?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ����?���Ǐ�?      �?        �q�q�?�8��8��?              �?      �?        ۬�ڬ��?�LɔL��?8��Moz�?d!Y�B�?�������?�������?              �?�m۶m��?�$I�$I�?              �?      �?        F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?        �׽�u��?�E(B�?�m۶m��?�$I�$I�?      �?      �?      �?        �������?�������?�$I�$I�?۶m۶m�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        ;�;��?��؉���?�������?ZZZZZZ�?      �?      �?���L�?}���g�?�������?""""""�?�������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?�������?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?      �?        �������?�������?      �?                      �?      �?              �?        O����?�}�+r��?|�)�C�?{>�e�ī?�a�a�?��y��y�?              �?�t�V�?9��v���?�?�?��8��8�?�q�q�?      �?        [4���?'u_[�?�7��Mo�?d!Y�B�?      �?        xxxxxx�?�?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �Y�	qV�?�cj`?      �?        �F��F��?�5�5�?��.���?t�E]t�?      �?        �������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �D�a�Y�?���Id�?Hy�G�?�n�ᆫ?.�u�y�?;ڼOqɐ?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?9��8���?�q�q�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?ӛ���7�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?۶m۶m�?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        �������?�������?      �?              �?      �?      �?        ��}A�?�}A_З?      �?        _�_��?�A�A�?      �?        �?�?              �?      �?        N6�d�M�?e�M6�d�?333333�?�������?�������?�?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?333333�?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?333333�?              �?      �?              �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMChvh)h,K ��h.��R�(KMC��h}�B�P         r                 `f�$@��t���?�           8�@                                    @z�G�z�?�            @p@        ������������������������       �                      @               k                   @@@Z���c��?�            �o@                                   �?�۲I <�?�            �j@                                �|Y=@T�7�s��?#            �L@                                ���@"pc�
�?             &@               	                   �2@�q�q�?             @        ������������������������       �                     �?        
                        �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                03@�LQ�1	�?             G@                               ���@���"͏�?            �B@                                   �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@                                   �?�q�q�?             8@                               ��@�LQ�1	�?             7@        ������������������������       �                      @                                   �?����X�?             5@                                  �?�q�q�?             2@        ������������������������       �                     @                                ���@؇���X�?	             ,@        ������������������������       �                     �?        ������������������������       �8�Z$���?             *@        ������������������������       �                     @        ������������������������       �                     �?                                   �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        !       4                    �?�IA��?e            �c@        "       3                 �|Y>@     ��?             0@       #       2                    �?���Q��?             .@       $       -                   �6@և���X�?             ,@       %       ,                 xF� @X�<ݚ�?             "@       &       +                    �?r�q��?             @       '       *                   �3@z�G�z�?             @        (       )                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        .       /                 �&B@z�G�z�?             @        ������������������������       �                      @        0       1                    9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        5       H                 �?�@`	�<��?V            �a@       6       E                   �?@��p\�?.            �T@       7       <                 ���@ �\���?,            �S@        8       9                    7@����X�?             @        ������������������������       �                     @        :       ;                 �&b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        =       D                 �?$@������?'             R@        >       ?                 �|Y;@HP�s��?             9@       ������������������������       �        
             2@        @       C                 �|Y>@����X�?             @       A       B                 ��@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �G@        F       G                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       R                 @3�@��$�4��?(            �M@        J       Q                    �?X�<ݚ�?             "@       K       P                    �?      �?              @       L       M                   �9@և���X�?             @        ������������������������       �                      @        N       O                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        S       h                 �|�=@j�q����?"             I@       T       a                 @�!@��0{9�?             �G@       U       ^                   � @"pc�
�?            �@@       V       ]                 0S5 @�>4և��?             <@       W       \                   �4@�+$�jP�?             ;@        X       Y                    1@X�<ݚ�?             "@        ������������������������       �      �?             @        Z       [                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     2@        ������������������������       �                     �?        _       `                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        b       c                 ���"@@4և���?
             ,@        ������������������������       �                     @        d       e                   �<@ףp=
�?             $@       ������������������������       �                     @        f       g                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        i       j                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        l       m                   @C@P�Lt�<�?             C@        ������������������������       �                     3@        n       o                    �?�}�+r��?             3@        ������������������������       �                      @        p       q                   �C@�IєX�?
             1@        ������������������������       ��q�q�?             @        ������������������������       �                     ,@        s                           @.iI\��?           0|@       t       �                  x#J@$;hB��?�            @s@       u       �                   �<@��U��?�            �j@        v       �                    �?��V#�?1            �U@       w       x                    �?@3����?             K@        ������������������������       �                      @        y       �                    �?��<b�ƥ?             G@        z       {                   �6@�nkK�?	             7@        ������������������������       �                     "@        |                          �9@@4և���?             ,@        }       ~                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     7@        �       �                    �?     ��?             @@        �       �                    �?և���X�?             @       �       �                   �8@���Q��?             @       �       �                 hf:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@HP�s��?             9@       ������������������������       �                     7@        ������������������������       �                      @        �       �                    �?b����?R            �_@       �       �                  �?@�8�Վ��?Q            @_@       �       �                    �?D��ٝ�?B            @Y@        �       �                    �?�eP*L��?             6@        �       �                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @C@     ��?	             0@       �       �                 ��";@r�q��?             (@       �       �                   @@@�q�q�?             @        ������������������������       �                     @        �       �                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���%&�?5            �S@       �       �                   �F@^H���+�?2            �R@       �       �                   @F@�[�IJ�?             �G@       �       �                   @E@�lg����?            �E@       �       �                     �?�e����?            �C@        �       �                 �|�?@�q�q�?             @       �       �                   �>@z�G�z�?             @       �       �                 `f�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �C@4���C�?            �@@       �       �                   @B@����"�?             =@       �       �                    �?
;&����?             7@        ������������������������       �                     "@        �       �                    1@؇���X�?             ,@       �       �                   �'@�<ݚ�?             "@        ������������������������       �                     @        �       �                    @@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �,@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �R@�<ݚ�?             ;@       �       �                    �?���B���?             :@        ������������������������       �                     @        �       �                    �?���}<S�?             7@       �       �                   �I@�C��2(�?             6@       �       �                 ��:@r�q��?             (@       ������������������������       �                      @        �       �                 `f�;@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             8@        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                     �?        �                         �O@�q�q�?A             X@       �       �                   �5@���!pc�?>             V@        �       �                   �1@��.k���?             1@       �       �                 ��f`@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 `fmj@@���?T�?3            �Q@       �       �                    �?     8�?.             P@       �       �                 ���P@���-T��?-             O@        �       �                 03sP@�z�G��?             4@       �       �                    �?@�0�!��?             1@        ������������������������       �                     $@        �       �                   �H@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                 0�nL@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?@4և���?              E@       �       �                    �?@-�_ .�?            �B@       �       �                    �?`Jj��?             ?@       ������������������������       �                     0@        �       �                    �?�r����?             .@        ������������������������       �                     @        �       �                   �H@      �?              @       �       �                 ЈT@؇���X�?             @        ������������������������       �                     @        �       �                   �D@      �?             @        ������������������������       �                      @        �       �                 Ј�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��W@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?և���X�?             @        ������������������������       �                     �?        �                          �?      �?             @                              �̾w@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                 �?x�f��^�?[            �a@                                 �?�>$�*��?            �D@                             X�,A@��+7��?             7@             	                  �0@��s����?             5@        ������������������������       �                     @        
                        �7@������?             .@        ������������������������       �                     �?                              �|Y=@d}h���?             ,@        ������������������������       �                      @                                 �?      �?             (@                              S�-@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             2@                             03�-@�eP*L��?             &@                                 3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r�q��?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              8                   �?t�F�}�?B            �Y@              /                   �?�q�q�?'             N@        !      *                ���5@*;L]n�?             >@       "      )                  �D@     ��?
             0@       #      (                   7@�r����?	             .@        $      '                   �?      �?             @       %      &                   +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        +      .                  @C@����X�?             ,@        ,      -                X��@@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0      1                   )@������?             >@        ������������������������       �                     @        2      7                   ;@H%u��?             9@        3      6                   �?և���X�?             @        4      5                �!&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        9      B                   @@4և���?             E@        :      ;                   �?���!pc�?             &@        ������������������������       �                     @        <      =                   @և���X�?             @        ������������������������       �                     @        >      ?                   �?      �?             @        ������������������������       �                      @        @      A                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �t�bh�h)h,K ��h.��R�(KMCKK��h^�B0  �nԾ���?5"W��6�?�������?�������?      �?        Y�eY�e�?��i��i�?T�rp�_�?��4>2��?p�}��?�}��?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?Nozӛ��?d!Y�B�?v�)�Y7�?*�Y7�"�?�؉�؉�?;�;��?              �?      �?        UUUUUU�?UUUUUU�?Nozӛ��?d!Y�B�?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        ;�;��?;�;��?      �?              �?        �q�q�?9��8���?              �?      �?        �(S�\��?�\�:�2�?      �?      �?333333�?�������?�$I�$I�?۶m۶m�?�q�q�?r�q��?UUUUUU�?�������?�������?�������?      �?      �?              �?      �?                      �?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?o����?E�)͋?�?�]�ڕ��?��+Q��?���7a�?�3���?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?q=
ףp�?{�G�z�?      �?        �m۶m��?�$I�$I�?333333�?�������?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        #h8����?u_[4�?r�q��?�q�q�?      �?      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?      �?              �?      �?        =
ףp=�?
ףp=
�?m�w6�;�?L� &W�?/�袋.�?F]t�E�?�$I�$I�?�m۶m��?/�����?B{	�%��?�q�q�?r�q��?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?              �?        �������?�������?      �?                      �?n۶m۶�?�$I�$I�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���k(�?(�����?      �?        �5��P�?(�����?      �?        �?�?UUUUUU�?UUUUUU�?      �?        �P�	e��?�^��5��?������?���8+?�?�[�琚�?tHM0���?6eMYS��?eMYS֔�?h/�����?���Kh�?              �?d!Y�B�?��7��M�?d!Y�B�?�Mozӛ�?              �?�$I�$I�?n۶m۶�?�������?�������?      �?                      �?              �?              �?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        q=
ףp�?{�G�z�?      �?                      �?5M�4M��?�eY�eY�?ˡE����?j�t��?�7���S�?z��~�X�?t�E]t�?]t�E�?UUUUUU�?�������?              �?      �?              �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        �g *��?�0���M�?L�Ϻ��?�g�`�|�?���
b�?m�w6�;�?}A_��?�}A_��?�-��-��?�A�A�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?                      �?m��&�l�?'�l��&�?	�=����?�i��F�?Y�B��?�Mozӛ�?              �?۶m۶m�?�$I�$I�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?      �?              �?      �?                      �?9��8���?�q�q�?��؉���?ى�؉��?              �?ӛ���7�?d!Y�B�?]t�E�?F]t�E�?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?                      �?�������?�������?      �?                      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?�������?�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�������?�������?      �?                      �?Zas �
�?�'�K=�?      �?     ��?�RJ)���?[k���Z�?333333�?ffffff�?�������?ZZZZZZ�?              �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?              �?      �?              �?              �?        �$I�$I�?n۶m۶�?к����?S�n0E�?�B!��?���{��?              �?�?�������?              �?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?�������?�������?              �?      �?              �?        �$I�$I�?۶m۶m�?      �?              �?      �?333333�?�������?      �?                      �?              �?      �?         2ܫ`��?��G�>��?�����?�18���?Y�B��?zӛ����?�a�a�?z��y���?              �?�?wwwwww�?      �?        ۶m۶m�?I�$I�$�?              �?      �?      �?333333�?ffffff�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?]t�E�?t�E]t�?�������?�������?              �?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        777777�?�������?�������?�������?�������?""""""�?      �?      �?�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        wwwwww�?�?              �?)\���(�?���Q��?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        n۶m۶�?�$I�$I�?F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@D         J                    �?�4�O��?�           8�@               5                    �?r�=���?~            �h@                                  �?T �����?[             c@                                   �?�i�y�?$            �O@                                  �?`Ӹ����?            �F@        ������������������������       �                     6@                                    @���}<S�?             7@        ������������������������       �                     @        	       
                 ���@�����H�?             2@        ������������������������       �                      @        ������������������������       �        
             0@        ������������������������       �        
             2@                                    �?��Hg���?7            �V@                                   �?և���X�?             5@                                  �?���Q��?             4@                               `f�A@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @                                  �5@      �?              @        ������������������������       �                      @                                  �H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                ���@�~t��?*            @Q@        ������������������������       �        
             2@               4                    �?��x_F-�?             �I@              3                 �|�=@j�q����?             I@              *                    �?      �?             B@              %                   �:@���y4F�?             3@                                 �&�)@�q�q�?             @        ������������������������       �                     �?        !       "                   �8@z�G�z�?             @        ������������������������       �                     @        #       $                 �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        &       )                   @@8�Z$���?             *@        '       (                 �|=@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        +       .                 �|Y=@�t����?
             1@        ,       -                  ��@      �?             @        ������������������������       �                      @        ������������������������       �                      @        /       2                    �?�θ�?             *@       0       1                  s�@�z�G��?             $@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     �?        6       C                    �?8�A�0��?#             F@       7       <                 �|Y=@�LQ�1	�?             7@       8       ;                 03�-@r�q��?
             (@        9       :                    &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        =       B                    �?�eP*L��?	             &@       >       ?                   @E@r�q��?             @        ������������������������       �                     @        @       A                 <3gH@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        D       I                     @؇���X�?             5@       E       H                 �̾w@�θ�?             *@       F       G                    )@�C��2(�?
             &@        ������������������������       �                     �?        ������������������������       �        	             $@        ������������������������       �                      @        ������������������������       �                      @        K       �                    �?D����?C           �@        L       m                    �?�BA����?f            `d@        M       l                   �J@�7�QJW�?/            �R@       N       [                     @v���a�?.            @R@       O       P                   �6@$�q-�?             J@        ������������������������       �        	             2@        Q       Z                   �*@�t����?             A@        R       S                   �'@�	j*D�?
             *@        ������������������������       �                      @        T       U                    :@���|���?             &@        ������������������������       �                      @        V       W                   �B@�<ݚ�?             "@       ������������������������       �                     @        X       Y                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        \       k                    @�q�q�?             5@       ]       j                 @�"@�z�G��?             4@       ^       i                 `��!@և���X�?
             ,@       _       b                 ���@�q�q�?	             (@        `       a                 �|Y:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        c       d                    4@և���X�?             @        ������������������������       �                      @        e       f                 @3�@z�G�z�?             @       ������������������������       �                     @        g       h                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        n       �                 �D�H@��7��?7             V@       o       �                    @�{r٣��?'            �P@       p       q                    @JJ����?            �G@        ������������������������       �                     @        r       �                    �?�D����?             E@       s       �                    @\�Uo��?             C@       t       u                   �6@և���X�?            �A@        ������������������������       �                     @        v       }                     @     ��?             @@        w       x                   �7@      �?             (@        ������������������������       �                      @        y       |                    �?ףp=
�?             $@       z       {                    D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~                        �|Y=@�z�G��?             4@        ������������������������       �                     @        �       �                    �?���Q��?             .@        �       �                 ��1@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 `fV6@�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��T?@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 pfv2@p�ݯ��?
             3@        ������������������������       �                     @        �       �                    �?$�q-�?             *@        ������������������������       �                      @        �       �                 ��T?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    #@�C��2(�?             6@        ������������������������       �                     �?        �       �                 ���P@���N8�?             5@        ������������������������       �                     $@        �       �                 X�,@@�C��2(�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                 ���d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?PN��T'�?�            �u@        �       �                   �>@�j�'�=�?*            �P@        �       �                   �<@r�q��?             8@        ������������������������       �                     @        �       �                   �Q@��Q��?             4@       �       �                   @E@�E��ӭ�?             2@       �       �                 03:@d}h���?
             ,@        ������������������������       �                      @        �       �                 03k:@      �?             @        ������������������������       �                     �?        �       �                 �|�?@���Q��?             @       �       �                 `fF<@      �?             @        ������������������������       �                      @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    K@      �?             @       �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�<@��s����?             E@        ������������������������       �                     @        �       �                    �?�ݜ�?            �C@       �       �                   �E@4?,R��?             B@       �       �                  x#J@�E��ӭ�?             2@       ������������������������       �                     "@        �       �                 �|Y>@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 `f�K@����X�?             @        �       �                 `�iJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             2@        ������������������������       �                     @        �       �                    '@�W�{�5�?�            �q@        �       �                     @��H�}�?             9@        ������������������������       �                     @        �       �                 ���A@      �?
             2@       �       �                    @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                 �?�@0Oex�I�?�            @p@        �       �                     @p� V�?=            �Y@        ������������������������       �                     @        �       �                    ?@@��8��?9             X@       �       �                   �8@@�z�G�?.             T@        �       �                    7@ ���J��?            �C@       ������������������������       �                     ?@        �       �                 `fF@      �?              @        �       �                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �       �                 �&B@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        �                          �?P��-�?h            �c@       �       �                     @0�I��8�?T             _@        �       �                    F@dP-���?!            �G@       �       �                   @D@������?            �B@       �       �                   �3@�#-���?            �A@       �       �                   �(@ȵHPS!�?             :@        �       �                   �5@$�q-�?             *@        �       �                    &@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�<@8�Z$���?
             *@        ������������������������       �                     @        �       �                   �A@�q�q�?             @       �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �      �?              @        ������������������������       �                     $@        �                         @@@؇���X�?3            @S@       �       
                �|Y>@���*�?&             N@       �                       �!&B@�t����?!            �I@       �       �                   �1@�8��8��?             H@        ������������������������       �                     $@        �       �                   �2@�KM�]�?             C@        ������������������������       �                     �?        �       �                 ��) @�L���?            �B@        ������������������������       �                     4@        �                       @3�!@@�0�!��?             1@        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?                               �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �<@@4և���?             ,@       ������������������������       �                     &@                              �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              	                   ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �?@X�<ݚ�?             "@        ������������������������       �                     @                              ��I @�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                    �@@        �t�bh�h)h,K ��h.��R�(KMKK��h^�B  �X�>�?2�N����?&���0�?m����g�?��G��G�?�\�\�?AA�?�������?l�l��??�>��?              �?d!Y�B�?ӛ���7�?              �?�q�q�?�q�q�?      �?                      �?              �?؂-؂-�?��I��I�?۶m۶m�?�$I�$I�?�������?333333�?�������?�������?              �?      �?              �?      �?      �?        UUUUUU�?�������?              �?      �?              �?        �s��\�?)�3J���?      �?        �������?�?=
ףp=�?
ףp=
�?      �?      �?6��P^C�?(������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?                      �?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �������?�������?      �?      �?      �?                      �?ى�؉��?�؉�؉�?ffffff�?333333�?      �?              �?      �?      �?              �?                      �?颋.���?/�袋.�?d!Y�B�?Nozӛ��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?t�E]t�?]t�E�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?ى�؉��?�؉�؉�?]t�E�?F]t�E�?              �?      �?                      �?      �?        &�%�%��?�K�K�K�?���+�j�?$���?0��b�/�?t�@�t�?�4iҤI�?ٲe˖-�?;�;��?�؉�؉�?              �?�?<<<<<<�?;�;��?vb'vb'�?              �?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?333333�?ffffff�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?              �?        ]t�E]�?�E]t��?��|��?|���?��
br�?x6�;��?              �?�0�0�?z��y���?�5��P^�?6��P^C�?�$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?ffffff�?333333�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?        9��8���?�q�q�?              �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        ^Cy�5�?Cy�5��?              �?�؉�؉�?;�;��?      �?        �������?�������?      �?                      �?F]t�E�?]t�E�?      �?        �a�a�?��y��y�?              �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?&���^B�?h/�����?�&�l���?m��&�l�?UUUUUU�?UUUUUU�?              �?�������?ffffff�?�q�q�?r�q��?I�$I�$�?۶m۶m�?      �?              �?      �?              �?333333�?�������?      �?      �?      �?              �?      �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?z��y���?�a�a�?              �?\��[���?�i�i�?�8��8��?r�q��?�q�q�?r�q��?      �?        �q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        �ĩ�sK�?Fڱa��?
ףp=
�?{�G�z�?              �?      �?      �?�������?�������?      �?                      �?      �?        �^�^��?�����?����`�?��,�?      �?        UUUUUU�?UUUUUU�?�������?�������?��-��-�?�A�A�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?                      �?6��(S��?R��fu�?!�B!�?��{���?�����F�?W�+�ɵ?��g�`��?к����?�A�A�?_�_�?��N��N�?�؉�؉�?�؉�؉�?;�;��?�������?UUUUUU�?              �?      �?              �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?              �?      �?      �?        ۶m۶m�?�$I�$I�?""""""�?wwwwww�?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?        �k(���?(�����?              �?}���g�?L�Ϻ��?      �?        ZZZZZZ�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?333333�?�������?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM%hvh)h,K ��h.��R�(KM%��h}�B@I         �                 `f~I@�t����?�           8�@              S                    �?�����2�?�           h�@                                ��@V���#�?~            �g@                                �|Y:@�IєX�?             1@       ������������������������       �                     &@                                �&�@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        	                            @�.�8�?q            �e@        
                        ���*@�L#���?/            �P@                                `f�)@      �?             8@                                  �J@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?                                  �B@"pc�
�?	             &@                                  :@�����H�?             "@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   E@ qP��B�?            �E@       ������������������������       �                     ?@                                    �?�8��8��?             (@        ������������������������       �                     @                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               &                    @�k��V��?B            �Z@                %                    �?؇���X�?             ,@       !       $                    @      �?              @        "       #                 ��0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        '       D                 03�1@�+Fi��?;             W@       (       =                 �?�-@�ݜ����?'            �M@       )       ,                 �̌@�&!��?            �E@        *       +                   �2@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        -       .                   �1@:ɨ��?            �@@        ������������������������       �                     @        /       <                    �?PN��T'�?             ;@       0       1                 `�X!@���y4F�?             3@        ������������������������       �                     @        2       7                   �9@����X�?	             ,@       3       6                    4@      �?              @        4       5                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        8       9                    �?      �?             @        ������������������������       �                     �?        :       ;                    A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        >       ?                   �0@      �?
             0@        ������������������������       �                     �?        @       C                   �;@��S�ۿ?	             .@        A       B                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        E       H                    @"pc�
�?            �@@       F       G                    �?�����?             5@        ������������������������       �                      @        ������������������������       �                     3@        I       J                 0C�7@�q�q�?             (@        ������������������������       �                     �?        K       L                    �?���!pc�?             &@        ������������������������       �                     @        M       N                    @      �?              @        ������������������������       �                      @        O       R                    @      �?             @       P       Q                   @C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        T       m                 �?�@б΅t�?           �x@        U       l                    �?�wY;��?X             a@       V       k                 �Yu@     x�?S             `@       W       b                    �?���F6��?B            �X@        X       Y                 ���@�ݜ�?            �C@        ������������������������       �        	             .@        Z       [                   �6@�q�q�?             8@        ������������������������       �                      @        \       ]                  ��@��2(&�?             6@        ������������������������       �                     "@        ^       _                 �|Y=@�θ�?	             *@        ������������������������       �                     �?        `       a                 X��A@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        c       d                    7@(;L]n�?)             N@        ������������������������       �                     3@        e       j                 ��L@������?            �D@       f       g                 ���@�(\����?             D@        ������������������������       �                     5@        h       i                 ���@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                      @        n       �                     �?|;�c� �?�            pp@        o       t                 �|�<@�q�q�?              H@        p       q                   �;@؇���X�?             @        ������������������������       �                      @        r       s                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        u       �                    �?���?            �D@       v       �                  �>@�d�����?             C@       w       �                    K@���Q��?             9@       x       �                   �G@���Q��?
             .@       y       ~                    �?���Q��?             $@        z       {                 `f&;@      �?             @        ������������������������       �                      @        |       }                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                 03k:@      �?             @        �       �                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���=@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @        �       �                    �?��ݼ��?�            �j@       �       �                     @�r����?W            �`@        �       �                    �? "��u�?              I@        ������������������������       �                     �?        �       �                    �?��<D�m�?            �H@       �       �                   �*@      �?             H@       �       �                 `fF)@l��\��?             A@        ������������������������       �                     $@        �       �                 �|�<@      �?             8@        ������������������������       �                     *@        �       �                   �F@���!pc�?             &@       �       �                 �|�=@      �?             @        ������������������������       �                     �?        �       �                    B@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     �?        �       �                    �?@�0�!��?7            @U@        ������������������������       �                     @        �       �                 @3�@����!�?4            �T@        �       �                    :@�eP*L��?             &@        ������������������������       �                     @        �       �                   �?@����X�?             @        ������������������������       �                      @        �       �                   �A@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        �       �                    )@D��\��?-            �Q@        ������������������������       �                     �?        �       �                 �|Y=@������?,            �Q@        �       �                 ��Y @��a�n`�?             ?@        �       �                   �3@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `�X#@�㙢�c�?             7@       �       �                 ���"@���y4F�?             3@       �       �                 @�!@�r����?
             .@       �       �                 pf� @�<ݚ�?             "@        ������������������������       �                      @        �       �                    8@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �?@�7��?            �C@       �       �                 ��) @���}<S�?             7@       ������������������������       �                     ,@        �       �                 �|�=@�<ݚ�?             "@       �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                    �?�z�G��?5             T@        �       �                 �2@�n_Y�K�?             *@       �       �                 �|�;@�����H�?             "@       �       �                 �&�)@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���}D�?-            �P@        �       �                    �? ��WV�?             :@        ������������������������       �                     @        �       �                    6@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    @��]�T��?            �D@       �       �                    �?\�Uo��?             C@        ������������������������       �                      @        �       �                    @�q�q�?             B@       �       �                 03{3@�q�����?             9@        �       �                     @z�G�z�?             $@        �       �                    *@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �̌4@�q�q�?             .@        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                    :@�z�G��?             $@       �       �                     @      �?             @        ������������������������       �                      @        �       �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                 pf�C@�q�q�?             @        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ƆQ����?P            �^@       �       �                  "�b@pY���D�?0            �S@       ������������������������       �        %            �M@        �       �                    �?ףp=
�?             4@       ������������������������       �                     $@        �       �                    $@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �                           @�&!��?             �E@       �                          �?p�ݯ��?             C@       �                           �?b�2�tk�?             B@       �       	                �UwR@���Q��?            �A@        �                          �?�<ݚ�?             2@                                  �?���Q��?             @        ������������������������       �                      @                              ��UO@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �C@$�q-�?             *@        ������������������������       �                     @                                 F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        
                         �?j���� �?             1@                                 �?      �?              @                                �?؇���X�?             @                                �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                                �?z�G�z�?             @                              �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @                                =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @              $                p�O@���Q��?             @              #                   >@      �?             @       !      "                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�b�d     h�h)h,K ��h.��R�(KM%KK��h^�BP  G�+J>�?r%�k���?37ı��?���w���?&N��[��?�X�0Ҏ�?�?�?              �?UUUUUU�?�������?      �?                      �?�avp��?+���}��?g��1��?��@���?      �?      �?;�;��?�؉�؉�?              �?      �?        F]t�E�?/�袋.�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?�}A_З?��}A�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?      �?                      �?����!5�?萚`���?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?              �?���,d!�?����7��?W'u_�?�}ylE��?֔5eMY�?S֔5eM�?333333�?ffffff�?      �?                      �?N6�d�M�?e�M6�d�?              �?&���^B�?h/�����?6��P^C�?(������?      �?        �m۶m��?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?        �������?333333�?              �?      �?              �?              �?      �?      �?        �?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?/�袋.�?F]t�E�?=��<���?�a�a�?              �?      �?        UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?      �?              �?      �?      �?              �?      �?�������?333333�?              �?      �?              �?        ��]�v��?�M�6%��?ZZZZZZ�?ZZZZZZ�?     @�?      �?�v�ļ�?ogH���?\��[���?�i�i�?      �?        UUUUUU�?�������?              �?��.���?t�E]t�?      �?        ى�؉��?�؉�؉�?              �?�������?UUUUUU�?�������?�������?      �?        �������?�?      �?        p>�cp�?������?333333�?�������?      �?        �5��P�?(�����?              �?      �?                      �?      �?              �?        ��4f��?���-g:�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        28��1�?8��18�?Cy�5��?y�5���?333333�?�������?�������?333333�?333333�?�������?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?      �?              �?      �?              �?                      �?�������?�������?      �?                      �?      �?              �?        =��˳��?��0�?�������?�?�G�z�?���Q��?      �?        ��S�r
�?և���X�?      �?      �?------�?�������?      �?              �?      �?      �?        F]t�E�?t�E]t�?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        ZZZZZZ�?�������?      �?        %jW�v%�?jW�v%j�?t�E]t�?]t�E�?      �?        �$I�$I�?�m۶m��?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?�o�z2~�?�@�6�?              �?,��+���?PuPu�?�c�1��?�s�9��?      �?      �?              �?      �?        �7��Mo�?d!Y�B�?6��P^C�?(������?�������?�?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?              �?      �?      �?                      �?      �?        ��[��[�?�A�A�?ӛ���7�?d!Y�B�?      �?        9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?        ffffff�?333333�?ى�؉��?;�;��?�q�q�?�q�q�?      �?      �?              �?      �?      �?      �?                      �?              �?      �?        &���[�?g��1��?O��N���?;�;��?      �?        �Mozӛ�?d!Y�B�?              �?      �?        KԮD�J�?jW�v%j�?�5��P^�?6��P^C�?      �?        �������?�������?���Q��?�p=
ף�?�������?�������?�������?�������?      �?                      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?ffffff�?333333�?      �?      �?              �?      �?      �?              �?      �?              �?                      �?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �}�K�`�?�`mާ�?�3���?a~W��0�?              �?�������?�������?              �?�������?�������?      �?                      �?֔5eMY�?S֔5eM�?^Cy�5�?Cy�5��?�8��8��?9��8���?333333�?�������?9��8���?�q�q�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ZZZZZZ�?�������?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        r�q��?�q�q�?�������?�������?      �?      �?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?      �?              �?        �������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK���h}�B�?                             @��ϙLq�?�           8�@               	                    @     ��?             @@                                  @��.k���?             1@                                  �?ףp=
�?             $@                                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        
                           �?��S�ۿ?
             .@       ������������������������       �                     $@                                   @z�G�z�?             @        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                 `fK@�ĸۦ��?�           8�@              Q                    �?��J��?r           @�@               "                     @Z�2�t��?h            �d@               !                    �?0)RH'�?(            @Q@                                 �*@�q�q��?             H@                                   B@���Q��?             4@                                 �9@      �?	             0@                                  �'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @                                ���;@ �Cc}�?             <@       ������������������������       �                     6@                                 X��C@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     5@        #       0                 pF @�W*��?@            @X@        $       /                    �?��hJ,�?             A@       %       .                 X��B@<���D�?            �@@       &       '                   �6@     ��?             @@        ������������������������       �                     .@        (       )                   �8@@�0�!��?             1@        ������������������������       �                      @        *       -                 ���@��S�ۿ?             .@        +       ,                 �Y�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     �?        ������������������������       �                     �?        1       N                 03�7@����X�?+            �O@       2       K                    �?�D����?             E@       3       F                    �?p�ݯ��?             C@       4       ?                 ��.@     ��?             @@       5       >                    �?�J�4�?             9@       6       ;                 �&�%@������?             1@       7       :                 `��!@ףp=
�?             $@        8       9                 `�X!@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        <       =                 ���*@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        @       A                    �?؇���X�?             @        ������������������������       �                     @        B       C                 03�1@      �?             @        ������������������������       �                      @        D       E                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        G       J                    @�q�q�?             @       H       I                   �4@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        L       M                 �|Y=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        O       P                    �?���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        R       �                   �J@T�1!�}�?
            z@       S       \                   �2@      �?�            �x@        T       [                 �&@������?             B@        U       V                    �?�X�<ݺ?             2@       ������������������������       �                     $@        W       Z                    �?      �?              @        X       Y                  �K"@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ]       x                     �?4�<����?�            @v@        ^       e                 �|�<@��J�fj�?            �B@        _       `                    7@      �?              @        ������������������������       �                     �?        a       b                 `f�D@؇���X�?             @       ������������������������       �                     @        c       d                 ��I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       w                   �G@J�8���?             =@       g       r                 �TA@@l��
I��?             ;@       h       m                 ���=@j���� �?             1@       i       l                 ��";@"pc�
�?
             &@       j       k                 ��:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        n       o                  �>@r�q��?             @        ������������������������       �                     @        p       q                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �C@ףp=
�?             $@       ������������������������       �                     @        u       v                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                    �?0�\>��?�            �s@       z       �                   @E@�u����?�             q@       {       �                    �?Ǖi�7�?�            0p@       |       �                     @X�EQ]N�?�             p@        }       ~                    �?���c���?             J@        ������������������������       �                     @               �                   @D@؇���X�?            �H@       �       �                 `fF)@�����H�?            �F@        �       �                    5@���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 �|�<@�㙢�c�?             7@        ������������������������       �                      @        �       �                   �3@������?             .@       �       �                   �A@�	j*D�?             *@       �       �                    @@      �?              @       �       �                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �      �?             @        �       �                 �Y�@�"�_*d�?�            �i@        �       �                   �8@���y4F�?             C@        �       �                   �3@���|���?             &@        ������������������������       �                     @        �       �                    5@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@ 7���B�?             ;@       ������������������������       �                     6@        ������������������������       �z�G�z�?             @        �       �                 �?�@4և����?k             e@       �       �                 �?$@x��B�R�?9            �V@        �       �                    ;@�8��8��?             B@        ������������������������       �                     *@        �       �                  s�@�LQ�1	�?             7@        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                 �|Y=@"pc�
�?	             &@        ������������������������       �                     �?        �       �                 X��A@ףp=
�?             $@       ������������������������       ������H�?             "@        ������������������������       �                     �?        �       �                 �|Y>@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                    �K@        �       �                    �?� ���?2            @S@        ������������������������       �                     @        �       �                   @C@�MI8d�?/            �R@       �       �                   �3@؇���X�?,            �Q@        ������������������������       ����Q��?             @        �       �                 ��) @�?�<��?*            @P@       �       �                   �>@��(\���?             D@       ������������������������       �                     =@        �       �                   �@@���!pc�?             &@       �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                     @        �       �                 �|�>@z�G�z�?             9@       �       �                   �8@      �?             4@        ������������������������       �                     @        �       �                 0S%"@     ��?             0@        �       �                 �|Y<@���Q��?             @        ������������������������       �                      @        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@"pc�
�?             &@        ������������������������       �                     @        �       �                 �|Y=@���Q��?             @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @D@      �?             @       �       �                 ��	0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 ��.@`Ӹ����?            �F@        �       �                    �?r�q��?	             (@       �       �                     @�C��2(�?             &@        ������������������������       �                     �?        �       �                    5@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     :@        �       �                    �?�"�q��?A            �W@       �       �                    �?�}�+r��?'            �L@       ������������������������       �                     =@        �       �                    @ �Cc}�?             <@       ������������������������       �                     9@        ������������������������       �                     @        �       �                    �?p�ݯ��?             C@       �       �                 X�,@@��Q��?             4@       �       �                  �}S@      �?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@       �       �                   @H@�����H�?             "@       ������������������������       �                     @        �       �                   �T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @b�2�tk�?             2@       �       �                     �?      �?	             (@       �       �                 �|Y>@�eP*L��?             &@        ������������������������       �                     �?        �       �                    �?���Q��?             $@       �       �                 03�U@      �?              @       �       �                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  �Ӭ����?�X�>��?      �?      �?�?�������?�������?�������?      �?      �?      �?                      �?              �?      �?        �?�������?              �?�������?�������?              �?      �?      �?      �?                      �?��T��?��W��?����Ǐ�?8p��?>�b���?፦ί=�?F��Q�g�?��k��?UUUUUU�?�������?�������?333333�?      �?      �?�������?�������?              �?      �?                      �?      �?        ۶m۶m�?%I�$I��?              �?      �?      �?              �?      �?                      �?�Q�/�~�?_\����?�������?KKKKKK�?|���?|���?      �?      �?              �?�������?ZZZZZZ�?      �?        �?�������?      �?      �?              �?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?�0�0�?z��y���?^Cy�5�?Cy�5��?      �?      �?�z�G��?{�G�z�?xxxxxx�?�?�������?�������?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?      �?      �?              �?      �?        ��y��y�?�a�a�?              �?      �?        �O���?�?��#s�?      �?      �?�q�q�?�q�q�?��8��8�?�q�q�?      �?              �?      �?�������?�������?      �?                      �?      �?              �?        �׽�u��?�E(B�?�"�u�)�?к����?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�rO#,��?|a���?Lh/����?h/�����?�������?ZZZZZZ�?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?              �?�]�b;��?�U�$��?<�H��?"��uy�?���K�?q�a�
��?w�qG�?qG�wĽ?;�;��?�;�;�?      �?        ۶m۶m�?�$I�$I�?�q�q�?�q�q�?�.�袋�?F]t�E�?              �?      �?        �7��Mo�?d!Y�B�?      �?        wwwwww�?�?vb'vb'�?;�;��?      �?      �?      �?      �?              �?      �?              �?      �?      �?              �?              �?      �?���[m�?���O ��?6��P^C�?(������?F]t�E�?]t�E]�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?	�%����?h/�����?      �?        �������?�������?I�$I�$�?�m۶m۶?�����?��?UUUUUU�?UUUUUU�?      �?        ��Moz��?Y�B��?      �?              �?      �?/�袋.�?F]t�E�?              �?�������?�������?�q�q�?�q�q�?      �?        �������?�������?      �?      �?      �?              �?        L�S�?��O����?      �?        ��L���?L�Ϻ��?۶m۶m�?�$I�$I�?333333�?�������?�����? �����?�������?333333�?      �?        F]t�E�?t�E]t�?      �?      �?              �?333333�?�������?      �?        �������?�������?      �?      �?      �?              �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        /�袋.�?F]t�E�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?        ?�>��?l�l��?�������?UUUUUU�?]t�E�?F]t�E�?      �?        �������?�������?              �?      �?                      �?      �?              �?        |n�S���?a�+F�?(�����?�5��P�?              �?۶m۶m�?%I�$I��?              �?      �?        Cy�5��?^Cy�5�?ffffff�?�������?      �?      �?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?�������?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        9��8���?�8��8��?      �?      �?]t�E�?t�E]t�?      �?        �������?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        UUUUUU�?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM5hvh)h,K ��h.��R�(KM5��h}�B@M         F                    �?�u����?�           8�@                                   �?sYi9��?O            `a@                                    @\#r��?"            �N@                                 �H@��<b�ƥ?             G@       ������������������������       �                     E@                                   J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        	                           �?�q�q�?
             .@       
                           �?X�Cc�?	             ,@                                �&�)@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                `�@1@����X�?             @                                  @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?               E                 �U�X@�θ�?-            �S@              D                  �	U@��R[s�?*            �Q@              C                    �?��ga�=�?(            �P@              <                 ��<J@�'�`d�?'            �P@              9                    �?&y�X���?#             M@              6                    �?r�����?             �J@              5                 p�i@@��k=.��?            �G@              2                   `A@�I�w�"�?             C@              1                 �|�=@"pc�
�?            �@@                                    �?d}h���?             <@                                0C�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        !       (                    ;@���B���?             :@        "       '                 ���@�8��8��?             (@       #       $                 ��y@؇���X�?             @        ������������������������       �                     �?        %       &                   �7@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        )       *                 �|Y=@����X�?	             ,@        ������������������������       �                     �?        +       ,                     @�θ�?             *@        ������������������������       �                     �?        -       0                   @@      �?             (@       .       /                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        3       4                      @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        7       8                 �&�)@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                ��k/@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =       B                 ���Q@      �?              @       >       A                    �?      �?             @       ?       @                    F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        G                          �?��s�ɝ�?t           ��@       H       �                    �?>4և���?"            |@       I       z                    �?������?�            �w@        J       g                   �9@z�G�z�?2            �R@        K       `                   �6@�û��|�?             7@       L       _                 8#B2@������?             1@       M       N                   �1@���|���?
             &@        ������������������������       �                     �?        O       X                   �4@���Q��?	             $@       P       Q                    �?      �?             @        ������������������������       �                     �?        R       W                    3@���Q��?             @       S       T                 P��@      �?             @        ������������������������       �                     �?        U       V                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                     @      �?             @        ������������������������       �                     �?        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ]       ^                 pF�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        a       b                     @r�q��?             @        ������������������������       �                     �?        c       f                    8@z�G�z�?             @       d       e                 @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        h       i                    �?ȵHPS!�?!             J@        ������������������������       �                     $@        j       w                     @؇���X�?             E@       k       n                 `f&'@ >�֕�?            �A@        l       m                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        o       p                     �?�g�y��?             ?@        ������������������������       �                     *@        q       r                   �B@�X�<ݺ?             2@       ������������������������       �                     "@        s       v                   �*@�����H�?             "@        t       u                    D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        x       y                 �|�;@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        {       �                 ��$:@�Qb��?�            �r@       |       �                   @@@������?�            0p@       }       �                   �>@$�3c�s�?v            �g@       ~       �                 @3�@��I�� �?o            `f@              �                 �|Y=@��<D�m�?;            �X@        �       �                 ��@      �?             D@       �       �                  ��@z�G�z�?             9@       �       �                    �?�C��2(�?             6@        ������������������������       �                     �?        �       �                    7@�����?             5@       ������������������������       �                     (@        �       �                 ���@�<ݚ�?             "@        �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        �       �                 �|�=@ _�@�Y�?             M@       �       �                     @@3����?             K@        ������������������������       �                     &@        �       �                 ��@ qP��B�?            �E@       ������������������������       �                     6@        �       �                 �Y5@���N8�?
             5@        ������������������������       �z�G�z�?             @        ������������������������       �                     0@        ������������������������       �                     @        �       �                   �3@�
��P�?4            @T@        �       �                   �2@�d�����?             3@       �       �                 ��Y @ףp=
�?             $@        �       �                    1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���$@X�<ݚ�?             "@       �       �                 0S5 @����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��a�n`�?(             O@        ������������������������       �                     �?        �       �                 ��) @\#r��?'            �N@        ������������������������       �                     6@        �       �                    :@8�Z$���?            �C@        ������������������������       �                     .@        �       �                     @      �?             8@        �       �                 �|Y<@�8��8��?             (@        ������������������������       �                     @        �       �                     �?؇���X�?             @        ������������������������       �                      @        �       �                 �|�=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 0S%"@�q�q�?             (@        �       �                 pf� @z�G�z�?             @        ������������������������       �                      @        �       �                 �|Y<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �&B@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �@      �?              @        ������������������������       �                     @        �       �                 �?�@���Q��?             @        ������������������������       �                     �?        �       �                 ��I @      �?             @       �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        �       �                   @E@�J�T�?-            �Q@       �       �                 �?�@�X�<ݺ?             B@        ������������������������       �        
             1@        �       �                 @3�@�KM�]�?             3@        ������������������������       ��q�q�?             @        �       �                   @D@      �?             0@       ������������������������       �                     ,@        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        �       �                     �?X��ʑ��?            �E@       �       �                 ��yC@j���� �?             A@       �       �                   �A@����X�?             <@       �       �                 �T!@@�q�q�?             8@       �       �                   �J@���!pc�?             6@       �       �                 `fF<@�t����?	             1@       �       �                 �|�?@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   @>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `fF<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ;@�<ݚ�?             "@        �       �                 ��?P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@DX�\��?3            �Q@        �       �                    �?��2(&�?             6@       �       �                     @     ��?             0@        �       �                    2@����X�?             @        ������������������������       �                     �?        �       �                     �?r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �!@�����H�?             "@        �       �                 ��Y@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?Rg��J��?%            �H@        �       �                   @C@���|���?             &@       �       �                    �?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �                           @      �?             C@       �                         @D@��}*_��?             ;@       �                           �?�<ݚ�?             2@       �                       �|Y=@r�q��?	             (@                               ���M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?ףp=
�?             $@       ������������������������       �                     @                              `f�K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �@@�q�q�?             @       	      
                  �<@z�G�z�?             @        ������������������������       �                     �?                                �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �?�q�q�?             "@                             �CdQ@      �?              @        ������������������������       �                     @                                 �?���Q��?             @        ������������������������       �                      @                              ��#[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?"pc�
�?             &@                              ���.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              (                    @�^�����?R             _@                                 �? i���t�?$            �H@       ������������������������       �                     C@               !                   �?�eP*L��?             &@        ������������������������       �                     �?        "      '                   �?���Q��?             $@       #      $                    �?X�<ݚ�?             "@        ������������������������       �                      @        %      &                   :@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        )      4                   �?��n�?.            �R@        *      +                  �7@���Q��?            �A@        ������������������������       �                     (@        ,      1                ��T?@���}<S�?             7@       -      0                   @@�}�+r��?             3@        .      /                �|Y>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        2      3                ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@        �t�bh�h)h,K ��h.��R�(KM5KK��h^�BP  ���|3�? ����?��]tc�?5	Q�E��?XG��).�?��:��?d!Y�B�?��7��M�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�m۶m��?%I�$I��?۶m۶m�?�$I�$I�?              �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?              �?ى�؉��?�؉�؉�?X|�W|��?PuPu�?��[���?�1���?6�d�M6�?'�l��&�?��FX��?�i��F�?Dj��V��?�V�9�&�?g���Q��?br1���?����k�?�5��P�?/�袋.�?F]t�E�?I�$I�$�?۶m۶m�?      �?      �?      �?                      �?��؉���?ى�؉��?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?              �?        �m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?              �?      �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?              �?        �������?333333�?              �?      �?              �?        �������?UUUUUU�?              �?      �?        �������?�������?              �?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?              �?      �?        ��y��3�?��*��?�m۶m[�?�$I�$I�?@2�խ �?��3T���?�������?�������?��,d!�?8��Moz�?�?xxxxxx�?F]t�E�?]t�E]�?              �?�������?333333�?      �?      �?              �?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�������?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �؉�؉�?��N��N�?              �?�$I�$I�?۶m۶m�?�A�A�?��+��+�?      �?      �?              �?      �?        �B!��?��{���?              �?�q�q�?��8��8�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?      �?        ـl@6 �?��M�&�?��P��?�{�ո�?1���\A�?x6�;��?��#���?Ck��P�?��S�r
�?և���X�?      �?      �?�������?�������?]t�E�?F]t�E�?      �?        =��<���?�a�a�?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        #,�4�r�?�{a���?���Kh�?h/�����?      �?        ��}A�?�}A_З?      �?        ��y��y�?�a�a�?�������?�������?      �?              �?        ������?��ӭ�a�?Cy�5��?y�5���?�������?�������?      �?      �?      �?                      �?      �?        r�q��?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?�s�9��?�c�1Ƹ?      �?        ��:��?XG��).�?      �?        ;�;��?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        �������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?�q�q�?r�q��?      �?              �?      �?              �?333333�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        (�K=�?��V؜?��8��8�?�q�q�?      �?        �k(���?(�����?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?              �?        ��}A�?�}A_�?ZZZZZZ�?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?�?<<<<<<�?;�;��?�؉�؉�?      �?                      �?      �?      �?      �?                      �?�������?�������?      �?                      �?      �?                      �?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        �]�����?�D+l$�?��.���?t�E]t�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?        ��S�r
�??4և���?F]t�E�?]t�E]�?333333�?ffffff�?              �?      �?              �?              �?      �?B{	�%��?_B{	�%�?�q�q�?9��8���?UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        !�B�?���{��?����X�?/�����?              �?]t�E�?t�E]t�?      �?        �������?333333�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?              �?      �?                      �?:m���?�K~���?333333�?�������?              �?ӛ���7�?d!Y�B�?�5��P�?(�����?�������?�������?      �?                      �?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK���h}�B@?         .                   �3@�L*�<�?�           8�@               +                    @b�L�4��?P            �`@                                  �?�Sb(�	�?A             [@                                   �?���.�6�?             G@        ������������������������       �        
             2@                                    @ �Cc}�?             <@       ������������������������       �                     2@               	                    @�z�G��?             $@        ������������������������       �                     @        
                           �?      �?             @                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                �?�@�g�y��?#             O@        ������������������������       �                     ,@                                   �?      �?             H@        ������������������������       �                      @                                    �?�LQ�1	�?             G@                                   �?և���X�?             <@                                   @      �?
             8@                                  �2@      �?             @        ������������������������       �                      @                                  �'@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                ��Y @      �?             2@                                  1@ףp=
�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        !       "                    �?�<ݚ�?             2@        ������������������������       �                      @        #       $                 03{3@      �?             0@        ������������������������       �                     $@        %       *                    �?�q�q�?             @       &       )                    �?���Q��?             @       '       (                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   -@$�q-�?             :@        ������������������������       �                      @        ������������������������       �                     8@        /       p                    �?B�����?_           �@        0       A                     @tHN�?q             f@       1       >                   @L@X'"7��?H             [@       2       3                    �?T��,��?D            @Y@        ������������������������       �                     A@        4       =                    �?�����?-            �P@       5       6                   �B@@4և���?             E@       ������������������������       �                     =@        7       8                   @C@�θ�?	             *@        ������������������������       �                     �?        9       :                     �?r�q��?             (@        ������������������������       �                     @        ;       <                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     9@        ?       @                   �L@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        B       m                    @\X��t�?)            @Q@       C       l                 03�:@p�EG/��?%            �O@       D       S                    �?d��0u��?"             N@        E       R                    �?������?             >@       F       Q                 ��.@l��
I��?             ;@       G       H                 �|Y=@X�<ݚ�?	             2@        ������������������������       �                     �?        I       N                    �?��.k���?             1@        J       M                    �?�<ݚ�?             "@       K       L                 X�x&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       P                 �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        T       k                   @B@��S���?             >@       U       f                    �?�5��?             ;@       V       ]                    �?      �?             4@       W       Z                 ��� @��
ц��?             *@       X       Y                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                 ���)@և���X�?             @        ������������������������       �                      @        `       e                 03�1@���Q��?             @       a       d                   �0@      �?             @       b       c                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        g       h                    �?؇���X�?             @        ������������������������       �                     @        i       j                 �|�:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       o                 ���4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        q       �                 ��D:@\���(\�?�             y@       r       �                    �?\2R}�?�            r@        s       ~                 �|Y=@�θV�?,            @Q@        t       }                    �?����X�?
             ,@       u       z                    �?�q�q�?             (@       v       w                   �8@�z�G��?             $@        ������������������������       �                     @        x       y                   @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        {       |                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               �                 �|�=@�1�`jg�?"            �K@       �       �                    �?Du9iH��?            �E@        �       �                    �?$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        �       �                   `3@��S�ۿ?             >@       �       �                 ���@h�����?             <@        ������������������������       �                     $@        �       �                   @'@�X�<ݺ?
             2@       ������������������������       �$�q-�?             *@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   @4@�2�~w�?�            �k@        �       �                 pf� @      �?             0@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �<@ =[y��?y            �i@        ������������������������       �        '            @P@        �       �                   �*@��X�-�?R            `a@       �       �                     @�#-���?@            @Z@        �       �                   �F@r�q��?             8@       �       �                   @D@���y4F�?             3@       �       �                 `fF)@r�q��?             2@       ������������������������       �                     $@        �       �                 �|�=@      �?              @        ������������������������       �                      @        �       �                    @@r�q��?             @        ������������������������       �                     @        �       �                   @B@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���"@xdQ�m��?/            @T@       �       �                 ��@ �\���?-            �S@        ������������������������       �                     7@        �       �                 ��L@@4և���?!             L@        �       �                 �|Y>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �@@`'�J�?            �I@       �       �                 ��) @`Jj��?             ?@       �       �                 @3�@h�����?             <@       �       �                 �?�@��S�ۿ?             .@       ������������������������       �                     $@        ������������������������       �z�G�z�?             @        ������������������������       �                     *@        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             4@        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        �       �                 p�w@�/e�U��?A            �[@       �       �                    �?� �W�??            �Z@       �       �                    �?X�Cc�?4             U@        �       �                 @�pX@
;&����?             7@       �       �                    �?b�2�tk�?             2@       �       �                 �|�;@�eP*L��?             &@        ������������������������       �                      @        �       �                 ��2>@�q�q�?             "@        ������������������������       �                      @        �       �                    C@؇���X�?             @       ������������������������       �                     @        �       �                 �D D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��`E@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    R@�ɞ`s�?%            �N@       �       �                 03k:@�c�Α�?$             M@        ������������������������       �                      @        �       �                 �!fK@      �?#             L@       �       �                     �?z�G�z�?             D@       �       �                    <@��G���?            �B@        ������������������������       �                     �?        �       �                   �F@r�q��?             B@       �       �                    �?�E��ӭ�?             2@       �       �                   `@@�n_Y�K�?
             *@        �       �                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @J@�X�<ݺ?
             2@        �       �                 `f�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                     @�n_Y�K�?	             *@       �       �                    C@�<ݚ�?             "@       �       �                 �|Y>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    >@      �?             @       �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?�nkK�?             7@       �       �                    �?�8��8��?             (@        �       �                 ��UO@؇���X�?             @        ������������������������       �                     @        �       �                   @D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �t�b�(     h�h)h,K ��h.��R�(KK�KK��h^�B�  KY� ��?iM���{�?���-�?v���?�Kh/���?�Kh/��?Y�B��?���7���?              �?۶m۶m�?%I�$I��?              �?333333�?ffffff�?              �?      �?      �?      �?      �?              �?      �?              �?        �B!��?��{���?      �?              �?      �?      �?        d!Y�B�?Nozӛ��?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?�������?�������?      �?      �?              �?      �?                      �?�q�q�?9��8���?      �?              �?      �?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?      �?                      �?              �?              �?�؉�؉�?;�;��?              �?      �?        bc ��?<9����?��5K�O�?�2���?B{	�%��?Lh/����?�F�tj�?�]?[��?              �?���@��?g��1��?�$I�$I�?n۶m۶�?              �?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?��Moz��?!Y�B�?Y�eY�e�?�4M�4M�?wwwwww�?DDDDDD�?�?wwwwww�?h/�����?Lh/����?�q�q�?r�q��?              �?�?�������?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?              �?              �?�������?�?/�����?h/�����?      �?      �?�؉�؉�?�;�;�?�m۶m��?�$I�$I�?              �?      �?        UUUUUU�?�������?      �?                      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?UUUUUU�?              �?      �?        �������?�������?B��_��?�M�]��?̵s���?�Q�g���?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?ffffff�?333333�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?      �?        A��)A�?�־a�?qG�w��?w�qGܱ?�؉�؉�?;�;��?      �?                      �?�������?�?�m۶m��?�$I�$I�?      �?        ��8��8�?�q�q�?�؉�؉�?;�;��?      �?              �?      �?      �?                      �?      �?        ־a��?A��)A�?      �?      �?      �?      �?      �?                      �?      �?        �������?�������?      �?        �.���?ݘ��V��?�A�A�?_�_�?�������?UUUUUU�?6��P^C�?(������?�������?UUUUUU�?      �?              �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �5?,R�?X�<ݚ�?���7a�?�3���?      �?        n۶m۶�?�$I�$I�?333333�?�������?              �?      �?        �������?�?���{��?�B!��?�m۶m��?�$I�$I�?�������?�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?              �?        �^����?�B�I .�?�#蝺�?9��/Ċ�?%I�$I��?�m۶m��?Y�B��?�Mozӛ�?9��8���?�8��8��?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?        mާ�d�?&C��6��?5�rO#,�?�{a���?              �?      �?      �?ffffff�?ffffff�?#�u�)��?v�)�Y7�?              �?�������?UUUUUU�?�q�q�?r�q��?;�;��?ى�؉��?UUUUUU�?�������?      �?                      �?      �?              �?        ��8��8�?�q�q�?      �?      �?              �?      �?              �?              �?              �?      �?;�;��?ى�؉��?9��8���?�q�q�?333333�?�������?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM)hvh)h,K ��h.��R�(KM)��h}�B@J         r                    �?]@f�
�?�           8�@               a                    �?��K�"�?�            �q@              &                 `f�$@�e�U��?�            �m@               %                    �?��H�}�?              I@              "                    �?(���@��?            �G@                               �̌@���� �?            �D@                               ���@�r����?             >@               	                 �|Y:@����X�?             @        ������������������������       �                     @        
                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?���}<S�?             7@       ������������������������       �        	             0@                                   4@����X�?             @        ������������������������       �                     �?                                �&B@r�q��?             @                                 �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  �2@���|���?             &@        ������������������������       �                     �?                                ��� @�z�G��?             $@                               @3�@r�q��?             @                                 �8@�q�q�?             @        ������������������������       �                     �?                                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                !                  SE"@      �?             @        ������������������������       �                      @        ������������������������       �                      @        #       $                   �3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        '       `                 �QD@X�E)9�?v            �g@       (       E                    �?�<�}���?K            @^@       )       D                    @�? Da�?(            �O@       *       +                    �?\#r��?&            �N@        ������������������������       �                     @        ,       5                 `f�)@ �Cc}�?#             L@        -       .                 pF%@`2U0*��?             9@        ������������������������       �                     *@        /       0                    +@�8��8��?             (@        ������������������������       �                     @        1       4                    �?r�q��?             @       2       3                 ��&@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        6       =                   �*@�חF�P�?             ?@        7       <                   �B@X�<ݚ�?             "@       8       ;                    �?����X�?             @       9       :                    <@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        >       ?                    �?���7�?             6@       ������������������������       �                     .@        @       C                    1@؇���X�?             @       A       B                    "@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        F       _                   �@@V�a�� �?#             M@       G       H                    �?F�t�K��?"            �L@        ������������������������       �        	             .@        I       J                   �9@0,Tg��?             E@        ������������������������       �                     ,@        K       T                     @��>4և�?             <@       L       M                    6@      �?             0@        ������������������������       �                      @        N       S                    :@؇���X�?
             ,@       O       P                   �8@�<ݚ�?             "@        ������������������������       �                     �?        Q       R                   �E@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        U       ^                 �̤=@�q�q�?             (@       V       ]                 `fV6@�z�G��?             $@       W       X                 �|�;@և���X�?             @        ������������������������       �                     @        Y       Z                 03�1@      �?             @        ������������������������       �                      @        [       \                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        +             Q@        b       q                    @v�2t5�?            �D@       c       d                    �?      �?             A@        ������������������������       �                     @        e       f                     @�f7�z�?             =@        ������������������������       �                     @        g       h                    @�q�q�?             8@        ������������������������       �                     @        i       n                    *@p�ݯ��?
             3@       j       k                    @�8��8��?             (@        ������������������������       �                     @        l       m                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        o       p                 ���4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        s       �                 ��D:@���<��?           �z@       t       y                    $@�%�P��?�            �t@        u       v                     @"pc�
�?             &@        ������������������������       �                     @        w       x                 ��|2@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        z       �                     @ E�+0+�?�            �s@        {       |                   �)@�(\����?1             T@        ������������������������       �                    �A@        }       �                 ��,@`Ӹ����?            �F@       ~                        �|�<@$�q-�?             :@        ������������������������       �                     ,@        �       �                 �|�=@r�q��?             (@        ������������������������       �                     �?        �       �                   �A@�C��2(�?             &@       �       �                    @@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     3@        �       �                    �?��5Վ3�?�            �m@        �       �                    �?^������?            �A@       �       �                    �?�c�Α�?             =@       �       �                 ���@      �?             8@        ������������������������       �                     @        �       �                   @@�q�q�?
             2@        �       �                   �5@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �|=@և���X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        �       �                 �|�;@�����H�?             "@        �       �                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �&�)@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��y&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@@ ��fί�?�            `i@       �       �                    �?3��e��?j            �d@       �       �                   �:@$s��O�?Z            �a@        �       �                   �2@�FVQ&�?,            �P@        �       �                   �1@      �?
             (@       �       �                   �0@�<ݚ�?             "@       �       �                 pf�@����X�?             @        ������������������������       �                      @        �       �                 pFD!@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@�q�q�?             @        ������������������������       �                     �?        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@3����?"             K@        ������������������������       �                      @        �       �                 ���@ pƵHP�?!             J@        �       �                    7@z�G�z�?             @        ������������������������       �                      @        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �G@        �       �                 ��) @��A��?.            �R@       �       �                 @3�@lGts��?$            �K@       �       �                   �>@(L���?            �E@       �       �                 �|Y=@     ��?             @@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��(@�>����?             ;@       �       �                 03�@      �?             0@        ������������������������       �                     @        ������������������������       �"pc�
�?             &@        ������������������������       �                     &@        �       �                   �?@���!pc�?             &@        �       �                 pff@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     (@        �       �                 ��)"@p�ݯ��?
             3@        �       �                 �|Y<@      �?              @        ������������������������       �                     @        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�C��2(�?             &@        ������������������������       �                      @        �       �                    (@�����H�?             "@        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? 7���B�?             ;@       ������������������������       �                     6@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        �                          �J@*Mp����?J            �Y@       �       �                 ��";@|jq��?<            �T@        �       �                 03k:@      �?              @        ������������������������       �                     �?        �       �                 �|�?@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                   �C@      �?             @        ������������������������       �                     �?        �       �                    H@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                   �;@L�qA��?5            �R@        �       �                    6@l��[B��?             =@       �       �                    �?�����?             3@       ������������������������       �                     "@        �       �                    @���Q��?             $@        ������������������������       �                     @        �       �                    @�q�q�?             @       �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �                           �?���j��?!             G@       �                         �I@P����?             C@       �                          �?<ݚ)�?             B@       �                         �H@����X�?            �A@                              p�w@     ��?             @@                                �?������?             >@                             `f�B@�GN�z�?             6@                               �A@�eP*L��?	             &@             	                   �?�q�q�?             "@                              �|�=@�q�q�?             @        ������������������������       �                     �?                                �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                        �>@r�q��?             @                               @=@�q�q�?             @        ������������������������       �                     �?                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                                 �?      �?              @                             `ށK@և���X�?             @        ������������������������       �                      @                                �G@���Q��?             @                                @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        !      (                   �?�}�+r��?             3@       "      #                   �?$�q-�?	             *@        ������������������������       �                     @        $      '                 )?@r�q��?             @        %      &                  �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM)KK��h^�B�  ߺ?9���?C����v�?|�W|�W�?����?=����Y�?�UP����?
ףp=
�?{�G�z�?R�٨�l�?W�+���?,Q��+�?jW�v%j�?�?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?ӛ���7�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E]�?F]t�E�?              �?ffffff�?333333�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        p����?��G'��?�C��2(�?�GN��?AA�?�������?XG��).�?��:��?              �?۶m۶m�?%I�$I��?{�G�z�?���Q��?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?�������?�������?      �?                      �?              �?��RJ)��?�Zk����?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        F]t�E�?�.�袋�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        a���{�?��{a�?:��,���?1��t��?              �?1�0��?�y��y��?              �?I�$I�$�?۶m۶m�?      �?      �?      �?        �$I�$I�?۶m۶m�?�q�q�?9��8���?              �?      �?      �?              �?      �?                      �?�������?�������?ffffff�?333333�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?                      �?��+Q��?�ڕ�]��?      �?      �?              �?O#,�4��?a���{�?              �?�������?�������?      �?        ^Cy�5�?Cy�5��?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        K�M�x[�?��Ȳ��?'^O��?����?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?              �?      �?        �k#֥��?��N�¹?333333�?�������?      �?        ?�>��?l�l��?�؉�؉�?;�;��?      �?        �������?UUUUUU�?              �?]t�E�?F]t�E�?�������?UUUUUU�?      �?              �?      �?      �?              �?        e�e��?�k"�k"�?uPuP�?_�_��?5�rO#,�?�{a���?      �?      �?      �?        UUUUUU�?UUUUUU�?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?      �?        �������?333333�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?����)�?xÏ���?6�'���?S&���?�A�A�?_�_��?>����?|���?      �?      �?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ���Kh�?h/�����?      �?        'vb'vb�?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��g�`�?�g�`�|�?�<%�S��?�־a�?⎸#��?w�qG��?      �?      �?�������?�������?              �?      �?        �Kh/��?h/�����?      �?      �?      �?        /�袋.�?F]t�E�?      �?        F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?        ^Cy�5�?Cy�5��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?        �q�q�?�q�q�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        	�%����?h/�����?      �?        �������?�������?              �?      �?              �?        �?�������?��ί=��?�b��7�?      �?      �?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?t�@��?�K~���?GX�i���?���=��?Q^Cy��?^Cy�5�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        �������?�������?              �?      �?        ozӛ���?!Y�B�?�P^Cy�?Q^Cy��?��8��8�?�8��8��?�m۶m��?�$I�$I�?      �?      �?wwwwww�?�?�袋.��?]t�E�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?      �?              �?      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?                      �?              �?      �?        �5��P�?(�����?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM'hvh)h,K ��h.��R�(KM'��h}�B�I                             @	dm#��?�           8�@                                   @     ��?              H@                               �-]@(;L]n�?             >@       ������������������������       �                     <@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               	                    �?�<ݚ�?
             2@        ������������������������       �                     $@        
                        ��T?@      �?              @        ������������������������       �                      @                                   @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               "                  @L@^ɼ���?�           ��@              W                    �?@\L5�T�?�           ؃@               4                     @l��TO��?H            @_@                                  �?�M���?(             Q@                                03�=@�X�<ݺ?             B@                                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     <@               )                 �D�G@     ��?             @@                                 �;@��.k���?             1@        ������������������������       �                     �?               (                     �?     ��?
             0@              '                    �?��
ц��?             *@              &                    C@�q�q�?             (@              %                   �A@�eP*L��?             &@              $                 ��2>@���Q��?             $@               #                 �ܵ<@      �?              @       !       "                 X�,@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        *       +                  �}S@������?
             .@        ������������������������       �                     @        ,       3                    �?      �?              @       -       2                    �?�q�q�?             @       .       1                    �?      �?             @       /       0                   �=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        5       N                    �?�MWl��?             �L@       6       9                    �?:	��ʵ�?            �F@        7       8                 `�@1@      �?              @       ������������������������       �                     @        ������������������������       �                      @        :       G                 �|Y=@�MI8d�?            �B@        ;       @                 ���@X�Cc�?             ,@        <       =                    5@���Q��?             @        ������������������������       �                     �?        >       ?                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        A       F                   �<@�<ݚ�?             "@       B       C                   �8@      �?              @        ������������������������       �                     @        D       E                   @;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        H       I                 ���@�nkK�?             7@        ������������������������       �                     @        J       M                 �|�=@      �?             0@       K       L                   @@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        O       V                 ���.@�q�q�?             (@       P       U                    �?      �?              @       Q       R                    �?r�q��?             @        ������������������������       �                     @        S       T                 �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X                       0�^I@Gq����?F           �@       Y       �                     @�"��c��?           P|@        Z       �                    �?z�7�Z�?\            @b@       [       t                 �|Y=@$��fF?�?L            @_@        \       a                    &@H�z�G�?             D@        ]       ^                    �?X�Cc�?             ,@        ������������������������       �                     @        _       `                   �7@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        b       k                   �;@�	j*D�?             :@       c       f                    �?�t����?             1@        d       e                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       h                    :@��S�ۿ?             .@       ������������������������       �        	             (@        i       j                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    �?�q�q�?             "@        ������������������������       �                     @        n       s                 `f�D@���Q��?             @       o       p                 `fF<@�q�q�?             @        ������������������������       �                     �?        q       r                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        u       �                   �*@ܻ�yX7�?1            @U@        v       }                   �>@��p\�?            �D@        w       x                    �?�r����?
             .@        ������������������������       �                     �?        y       |                 �|�=@@4և���?	             ,@       z       {                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ~                           �? ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �2@���|���?             F@        ������������������������       �                     @        �       �                   @J@�z�G��?             D@       �       �                    �?�q�q�?             B@       �       �                    �?`�Q��?             9@        ������������������������       �                      @        �       �                     �?��+7��?             7@       �       �                   �>@�z�G��?             4@       �       �                 ��<:@�eP*L��?             &@        ������������������������       �                      @        �       �                 X��B@�q�q�?             "@        ������������������������       �                      @        �       �                    H@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?���|���?             &@        �       �                   �E@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    *@���N8�?             5@        ������������������������       �                      @        �       �                    �?�S����?             3@       ������������������������       �                     0@        ������������������������       �                     @        �       �                    �?4����?�            0s@        �       �                    �?      �?             L@        �       �                    @���B���?             :@       �       �                    �?���}<S�?             7@       �       �                 �|�9@      �?	             0@        ������������������������       �                     @        �       �                  ��@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     >@        �       �                    �?���w;�?�            `o@        �       �                    �?�G�5��?)            @Q@       �       �                 ���1@b�2�tk�?             B@       �       �                 �|�<@��S���?             >@       �       �                 pf�@�q�q�?             2@        ������������������������       �                     @        �       �                   �2@z�G�z�?	             .@        ������������������������       �                     @        �       �                    �?      �?             (@       �       �                   �@�<ݚ�?             "@        �       �                 �&B@�q�q�?             @       �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?	             (@        �       �                   &@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��Y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    :@�C��2(�?            �@@       �       �                   �6@@�0�!��?
             1@       �       �                   �0@��S�ۿ?	             .@       ������������������������       �                     "@        �       �                    3@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     0@        �       �                 �?�@|)����?z            �f@        �       �                    ?@@�)�n�?9            @U@       �       �                    �?�\=lf�?-            �P@       �       �                 ���@ ������?)            �O@        �       �                   �8@�����H�?             "@        �       �                   �4@z�G�z�?             @        ������������������������       �                     �?        �       �                 �&b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        #             K@        ������������������������       �                     @        �       �                 �&B@�����H�?             2@       ������������������������       �                     (@        �       �                   �A@�q�q�?             @        �       �                   �@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                          �?�*v��?A            @X@       �       �                 @3�@ ��~���?<            �V@        �       �                    �?X�Cc�?             ,@       �       �                   �A@�	j*D�?             *@       �       �                   �:@"pc�
�?             &@        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    )@�KM�]�?4             S@        ������������������������       �                     �?        �                          ?@���Lͩ�?3            �R@       �                       �|�=@H�ՠ&��?$             K@       �                          �?���C��?#            �J@       �                          �?�t����?!            �I@       �                       @3�!@(L���?            �E@       �       �                 �|Y<@@�0�!��?             A@       �       �                 pf� @      �?             0@       �       �                 0S5 @"pc�
�?	             &@       �       �                   �3@�<ݚ�?             "@        �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    8@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ��) @�����H�?
             2@       ������������������������       �                     .@        �                        pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @                                  @�q�q�?*            �L@       	      
                   �?���3�E�?%             J@       ������������������������       �                     @@                                 �?      �?             4@                                 �?�E��ӭ�?             2@                               �E@     ��?             0@                              x#J@�n_Y�K�?             *@        ������������������������       �                     @                                 �?      �?             $@        ������������������������       �                     �?                              `�iJ@X�<ݚ�?             "@        ������������������������       �                     @                              `f�N@�q�q�?             @                                7@      �?             @        ������������������������       �                     �?                                 A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @              !                   �?z�G�z�?             @                                  ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #      &                   �?h�����?             <@        $      %                  pE@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �t�bh�h)h,K ��h.��R�(KM'KK��h^�Bp  �"iD��?&�-w���?      �?      �?�?�������?              �?      �?      �?              �?      �?        9��8���?�q�q�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��Е���?�6^�6^�?[�V��j�?K�R�T*�?h��|?5�?L7�A`��?<<<<<<�?�������?�q�q�?��8��8�?      �?      �?      �?                      �?              �?      �?      �?�������?�?              �?      �?      �?�؉�؉�?�;�;�?�������?�������?]t�E�?t�E]t�?�������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?                      �?      �?              �?        �?wwwwww�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?:��,���?�YLg1�?��O��O�?l�l��?      �?      �?      �?                      �?��L���?L�Ϻ��?%I�$I��?�m۶m��?�������?333333�?      �?              �?      �?              �?      �?        9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�Mozӛ�?d!Y�B�?      �?              �?      �?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?        �������?�������?      �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?�������?�?o���?E�w<���?�I�&M��?�lٲe��?bX9���?;�O��n�?ffffff�?333333�?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?        vb'vb'�?;�;��?<<<<<<�?�?      �?      �?              �?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        �������?�������?�]�ڕ��?��+Q��?�������?�?              �?n۶m۶�?�$I�$I�?]t�E�?F]t�E�?      �?                      �?      �?        O��N���?;�;��?              �?      �?        ]t�E]�?F]t�E�?              �?ffffff�?333333�?UUUUUU�?UUUUUU�?��(\���?{�G�z�?              �?zӛ����?Y�B��?ffffff�?333333�?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��y��y�?�a�a�?      �?        ^Cy�5�?(������?              �?      �?        9T��_�?�����?      �?      �?ى�؉��?��؉���?d!Y�B�?ӛ���7�?      �?      �?              �?�������?�������?      �?                      �?              �?      �?              �?        ������?�핷$��?��v`��?�%~F��?�8��8��?9��8���?�?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?                      �?      �?        ]t�E�?F]t�E�?ZZZZZZ�?�������?�������?�?      �?        �������?UUUUUU�?              �?      �?                      �?      �?        ��/��/�?h�h��?�������?�?"=P9���?g��1��?��}��}�?AA�?�q�q�?�q�q�?�������?�������?      �?              �?      �?      �?                      �?      �?              �?              �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ��Id��?�i�n�'�?�`�`�?�'}�'}�?%I�$I��?�m۶m��?vb'vb'�?;�;��?/�袋.�?F]t�E�?      �?        333333�?�������?              �?              �?�k(���?(�����?              �?�6�i�?�K~��?������?{	�%���?\�琚`�?"5�x+��?<<<<<<�?�?⎸#��?w�qG��?ZZZZZZ�?�������?      �?      �?/�袋.�?F]t�E�?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        333333�?�������?      �?                      �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?                      �?      �?              �?        UUUUUU�?UUUUUU�?b'vb'v�?O��N���?              �?      �?      �?�q�q�?r�q��?      �?      �?;�;��?ى�؉��?      �?              �?      �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?              �?        �������?�������?      �?      �?              �?      �?              �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�C         P                     �?e�L��?�           8�@               3                    �?�G�z�?f             d@                                  �?���r
��?A            @X@                                   �?�D����?             E@                                 @H@p�ݯ��?             C@                               �|�;@�������?             >@        ������������������������       �                     &@               	                    �?p�ݯ��?             3@       ������������������������       �                     $@        
                          �A@�<ݚ�?             "@                               X�,@@����X�?             @                               ��2>@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                ��Z@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               *                 0�_J@N{�T6�?$            �K@                                  �?��.k���?             A@        ������������������������       �                     @                                �|�<@���Q��?             >@        ������������������������       �                     @               )                    R@�q�q�?             ;@              (                    L@�	j*D�?             :@              '                   �>@���Q��?             4@                                �̌*@�q�q�?             (@        ������������������������       �                      @        !       "                   �C@z�G�z�?             $@        ������������������������       �                     @        #       &                 `f�;@�q�q�?             @       $       %                    H@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        +       0                 03c@؇���X�?             5@       ,       -                    �?�IєX�?	             1@       ������������������������       �                     .@        .       /                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                 ���f@      �?             @        ������������������������       �                      @        ������������������������       �                      @        4       O                   �P@�<ݚ�?%            �O@       5       @                 ��Q@���*�?$             N@        6       7                    �?�q�q�?             2@        ������������������������       �                     @        8       ?                    F@�eP*L��?             &@       9       :                    �?r�q��?             @        ������������������������       �                      @        ;       >                   @B@      �?             @       <       =                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        A       H                    �?���H��?             E@       B       G                    �?`Jj��?             ?@       C       D                    �?$�q-�?             :@       ������������������������       �        
             2@        E       F                 ���^@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        I       L                    �?���!pc�?             &@       J       K                 �U�X@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        M       N                 ��f`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Q       �                    �?�w�+`�?]           8�@       R       �                 Ь�#@�;�T<:�?           �z@       S       T                 ���@D�a�ў�?�            �p@        ������������������������       �                     <@        U       V                 ��@�.�PI�?�            �m@        ������������������������       �                     @        W       X                    /@P�z�?�            `m@        ������������������������       �                      @        Y       p                    �?F�|���?�             m@        Z       [                    �?Dc}h��?&             L@        ������������������������       �        	             *@        \       i                    �?�ʈD��?            �E@       ]       h                 �� @�LQ�1	�?             7@       ^       a                 ���@؇���X�?             5@        _       `                 �|�9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        b       g                 �|Y=@r�q��?	             (@        c       d                   @8@�q�q�?             @        ������������������������       �                     �?        e       f                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        j       k                 ���@P���Q�?             4@        ������������������������       �                     @        l       o                 X�I@      �?             0@       m       n                 ��(@��S�ۿ?             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        ������������������������       �                     �?        q       v                    �?$���?f             f@        r       u                   �@
;&����?             7@        s       t                   �A@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     &@        w       �                 �?�@�C��2(�?Z            @c@       x       y                 �|�<@����D��?5            @W@       ������������������������       �                     J@        z       �                   @@@������?            �D@       {       �                   �@�8��8��?             8@        |       �                 �&B@����X�?             @       }       ~                 ��@r�q��?             @        ������������������������       �                     @               �                 �|Y>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     1@        �       �                   �4@`��:�?%            �N@        �       �                   �0@�q�q�?
             .@        ������������������������       ����Q��?             @        �       �                 @3�@�z�G��?             $@        ������������������������       �                      @        �       �                 ��Y @      �?              @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@*
;&���?             G@        �       �                   �A@      �?              @        ������������������������       �      �?             @        ������������������������       �      �?              @        �       �                    �?�˹�m��?             C@       �       �                 �|Y=@�8��8��?             B@        ������������������������       �                     "@        �       �                 �|Y?@�����H�?             ;@       �       �                 ��) @r�q��?	             2@       ������������������������       �                     &@        �       �                 pf� @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �       �                   �F@v�_���?e            �c@       �       �                   P,@�S��<�?Y            �a@        �       �                    �?      �?$             N@        �       �                     @ 7���B�?             ;@       ������������������������       �                     4@        �       �                    �?؇���X�?             @       �       �                 �[$@r�q��?             @        ������������������������       �                     @        �       �                 ��&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �%@<���D�?            �@@        ������������������������       �                     @        �       �                     @8�Z$���?             :@       �       �                 �|�<@�8��8��?             8@       ������������������������       �                     &@        �       �                 �|�=@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        �       �                 pf�/@d�� z�?5            @T@        �       �                    1@      �?             0@        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                     @�4��?)            @P@       �       �                    �?؀�:M�?            �B@        �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   �;@����X�?             @        ������������������������       �                     �?        �       �                   �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 ���1@����X�?             <@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?R���Q�?             4@        �       �                   �2@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �.@�IєX�?             1@       ������������������������       �        	             ,@        �       �                    5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @X9����?U            �_@        �       �                   �6@�������?             A@        ������������������������       �        
             .@        �       �                 ��J@�\��N��?             3@       �       �                    @���Q��?             .@       �       �                    �?X�Cc�?             ,@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?R�(��?=            @W@        �       �                 X��B@���y4F�?             3@       �       �                    @r�q��?             2@       �       �                    �?d}h���?             ,@       �       �                    3@r�q��?	             (@       �       �                    &@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                       �̼6@^��4m�?0            �R@        �                       �̌5@�'�=z��?            �@@       �       �                   �*@*;L]n�?             >@        �       �                    (@�z�G��?             $@       ������������������������       �                     @        �       �                 xFT$@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�z�G��?             4@       �       �                     @8�Z$���?	             *@       �       �                    )@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                 @33/@և���X�?             @        ������������������������       �                     �?        �                           �?�q�q�?             @        ������������������������       �                     @                                 +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              
                   �?��p\�?            �D@              	                  @C@�t����?
             1@                                �B@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@                              ��p@@ �q�q�?             8@                              ��T?@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        
             *@        �t�b��     h�h)h,K ��h.��R�(KMKK��h^�B�  v�S(��?��X��?�������?�������?���fy�?�<�L�v�?z��y���?�0�0�?Cy�5��?^Cy�5�?�������?�������?              �?Cy�5��?^Cy�5�?              �?9��8���?�q�q�?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        pX���o�?�S�<%��?�������?�?              �?333333�?�������?              �?UUUUUU�?UUUUUU�?vb'vb'�?;�;��?333333�?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?              �?                      �?�$I�$I�?۶m۶m�?�?�?              �?      �?      �?              �?      �?              �?      �?      �?                      �?�q�q�?9��8���?wwwwww�?""""""�?UUUUUU�?UUUUUU�?              �?t�E]t�?]t�E�?UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��y��y�?�0�0�?�B!��?���{��?;�;��?�؉�؉�?              �?      �?      �?              �?      �?                      �?t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?      �?                      �?      �?        n�x�2��?%g����?\�琚`�?��`��}�?��"��X�?�iu�՝�?      �?        �@��@��?��F��F�?              �?N(��-�?�^��H��?              �?��љT;�?m�����?�$I�$I�?۶m۶m�?              �?A_���?�}A_з?��Moz��?Y�B��?۶m۶m�?�$I�$I�?�q�q�?�q�q�?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        ffffff�?�������?      �?              �?      �?�������?�?�؉�؉�?;�;��?      �?              �?        ($�z�?^o�?�?Y�B��?�Mozӛ�?UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E�?F]t�E�?P?���O�?X`��?      �?        p>�cp�?������?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        *.�u��?XG��).�?UUUUUU�?UUUUUU�?333333�?�������?ffffff�?333333�?              �?      �?      �?      �?      �?              �?      �?              �?        ���,d!�?8��Moz�?      �?      �?      �?      �?      �?      �?��P^Cy�?^Cy�5�?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?�������?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?              �?         *�3�?���M���?P$�Ҽ��?`��Z��?      �?      �?h/�����?	�%����?              �?�$I�$I�?۶m۶m�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?|���?|���?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?        ;�;��?;�;��?              �?      �?                      �?��"e���?x�5?,�?      �?      �?      �?      �?      �?                      �?      �?        �R+�R+�?�Z��Z��?E>�S��?v�)�Y7�?      �?      �?              �?�������?�������?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?              �?        �m۶m��?�$I�$I�?      �?      �?              �?      �?        333333�?333333�?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        I$�D"�?o���v��?�������?�������?              �?�5��P�?y�5���?333333�?�������?%I�$I��?�m۶m��?              �?      �?                      �?              �?M4�DM�?f�]v�e�?(������?6��P^C�?UUUUUU�?�������?۶m۶m�?I�$I�$�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?      �?        �|����?�S�n�?|��|�?|���?""""""�?�������?333333�?ffffff�?              �?333333�?�������?      �?                      �?ffffff�?333333�?;�;��?;�;��?/�袋.�?F]t�E�?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�]�ڕ��?��+Q��?<<<<<<�?�?      �?      �?      �?                      �?      �?        �������?UUUUUU�?]t�E�?F]t�E�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@A         d                    �?e�L��?�           8�@               _                    @<�T]���?�            �o@              \                    @Q��"�?�            `m@              G                 �|�=@��^���?�             m@                                  !@ܱ#_��?\            `b@        ������������������������       �                     ,@                                   '@���c�?T            �`@        ������������������������       �                     @        	                            @:�����?R            �_@        
                           �?���J��?"            �I@        ������������������������       �                     4@                                   �?�g�y��?             ?@                                  9@P���Q�?             4@                                   �?      �?             @                                 �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     &@               :                    �?���=A�?0             S@              %                 @� @     ��?)             P@                                 �6@��s����?             E@        ������������������������       �        
             4@                                  �9@���|���?             6@                                pf�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   ;@�E��ӭ�?             2@        ������������������������       �                      @               $                    �?     ��?             0@               #                 ���@d}h���?	             ,@        !       "                 �Y�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        &       1                    �?8�A�0��?             6@        '       (                   �,@      �?             (@        ������������������������       �                      @        )       0                    �?�z�G��?             $@       *       /                  S�-@�q�q�?             "@       +       .                 �|Y6@���Q��?             @       ,       -                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        2       9                 �|�:@���Q��?	             $@       3       8                    �?؇���X�?             @       4       5                  �#@      �?             @        ������������������������       �                      @        6       7                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ;       @                   �6@�q�q�?             (@        <       ?                   �3@z�G�z�?             @       =       >                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        A       B                 �|�:@և���X�?             @        ������������������������       �                      @        C       D                    �?z�G�z�?             @        ������������������������       �                      @        E       F                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        H       W                    �?�̨�`<�?8            @U@       I       J                   @B@؇���X�?%             L@       ������������������������       �                     ;@        K       V                 83'E@�c�Α�?             =@       L       O                     �?      �?	             0@        M       N                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       U                   �+@�<ݚ�?             "@       Q       T                     @�q�q�?             @       R       S                    D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        X       Y                     @XB���?             =@       ������������������������       �                     7@        Z       [                    C@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ]       ^                 ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        `       a                      @�t����?             1@        ������������������������       �                     @        b       c                 �|Y?@$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        e       �                 ��K.@�#2����?"           �|@       f       w                    �?�]l*7��?�            0r@        g       h                   �6@>���Rp�?             M@        ������������������������       �                     "@        i       n                 �|Y=@ i���t�?            �H@        j       m                    �?      �?             (@       k       l                   �<@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        o       p                 ���@@-�_ .�?            �B@        ������������������������       �                     .@        q       r                     @�C��2(�?             6@        ������������������������       �                     @        s       v                 �|�=@�����H�?	             2@       t       u                   @@"pc�
�?             &@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     @        x       �                    �?`�q��־?�             m@       y       �                 ���"@ �Cc��?�             l@       z       �                 ��@�1��?o            �e@        {       |                     @��v$���?*            �N@        ������������������������       �                     $@        }       �                 ���@���J��?#            �I@        ~                        ���@�IєX�?
             1@       ������������������������       �        	             0@        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�h����?E             \@       �       �                   �3@ ѯ��?B            �Z@        �       �                   �1@��2(&�?             6@        ������������������������       �                     &@        �       �                 �?�@���!pc�?             &@        ������������������������       �                     @        �       �                 ��Y @���Q��?             @       �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     �?        �       �                 �|Y=@@�)�n�?6            @U@        ������������������������       �                    �B@        �       �                   @@@      �?             H@       �       �                    ?@�#-���?            �A@       �       �                 �|�=@@4և���?             <@       �       �                  sW@HP�s��?             9@        ������������������������       �      �?             @        ������������������������       �                     5@        ������������������������       �                     @        �       �                 P�@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @        �       �                   @B@�t����?$            �I@       �       �                   �@@R���Q�?             D@       �       �                     @�ݜ�?            �C@       �       �                    5@���7�?             6@        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     1@        �       �                 `�X#@������?             1@       �       �                   �<@�	j*D�?             *@        ������������������������       �                     @        �       �                 �|Y=@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �|�=@����X�?             @        ������������������������       �                     @        �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@      �?l             e@       �       �                   @A@�Sb(�	�?D             [@       �       �                 `�/@�Y|���?A            �Y@        ������������������������       �                     @        �       �                    @�D��??            �X@       �       �                    �?^H���+�?3            �R@       �       �                    �?�Gi����?            �B@       �       �                    �?���|���?            �@@        �       �                      @�q�q�?             "@       �       �                 �|Y<@����X�?             @        �       �                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �?@      �?             8@       �       �                 `f�D@����X�?             5@       �       �                     �?��
ц��?	             *@       �       �                   �<@�q�q�?             "@        ������������������������       �                      @        �       �                 `fF<@և���X�?             @        ������������������������       �                      @        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 h"_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?V������?            �B@        �       �                    �?�<ݚ�?             "@       �       �                    ;@      �?              @       �       �                    �?���Q��?             @       �       �                 8�T@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    )@��X��?             <@        ������������������������       �                     @        �       �                 `fFJ@�����?             5@       ������������������������       �        
             .@        �       �                     �?�q�q�?             @       �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        �       �                     �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?�?�P�a�?(             N@       �       �                    H@r�q��?             E@       �       �                    �?`2U0*��?             9@       �       �                    �?      �?	             0@        ������������������������       �                     �?        �       �                   �F@��S�ۿ?             .@        �       �                 `fF:@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     "@        �                       �5L@ҳ�wY;�?             1@       �                        i?@������?
             .@       �       �                 `fF:@���|���?             &@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?                                  L@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �t�bh�h)h,K ��h.��R�(KMKK��h^�BP  v�S(��?��X��?�������?AA�?*Kq��k�?5���	%�?X�i���?j��FX�?���+��?B����?              �?�����?Є?�L�?      �?        �F��h4�?].���r�?�?______�?              �?�B!��?��{���?�������?ffffff�?      �?      �?      �?      �?              �?      �?                      �?              �?              �?�P^Cy�?��P^Cy�?      �?     ��?�a�a�?z��y���?              �?F]t�E�?]t�E]�?      �?      �?              �?      �?        r�q��?�q�q�?              �?      �?      �?۶m۶m�?I�$I�$�?333333�?�������?              �?      �?                      �?      �?        /�袋.�?颋.���?      �?      �?              �?333333�?ffffff�?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?333333�?�������?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?�$I�$I�?۶m۶m�?              �?�{a���?5�rO#,�?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?      �?              �?                      �?�{a���?GX�i���?              �?UUUUUU�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?�؉�؉�?;�;��?      �?                      �?F)b���?�Zw>���?ݷ�x���?A�;��?�i��F�?GX�i���?              �?/�����?����X�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        S�n0E�?к����?      �?        ]t�E�?F]t�E�?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?�m۶m��?�$I�$I�?      �?              �?        ��6���?r؃H{�?I�$I�$�?n۶m۶�?��#���?+���}��?.�u�y�?;ڼOqɐ?      �?        ______�?�?�?�?      �?                      �?      �?        �$I�$I�?۶m۶m�?n���4�?�@�Ե�?��.���?t�E]t�?      �?        F]t�E�?t�E]t�?      �?        �������?333333�?      �?      �?              �?      �?      �?      �?        �������?�?      �?              �?      �?�A�A�?_�_�?n۶m۶�?�$I�$I�?q=
ףp�?{�G�z�?      �?      �?      �?              �?        ۶m۶m�?�$I�$I�?              �?      �?              �?              �?        <<<<<<�?�?333333�?333333�?\��[���?�i�i�?�.�袋�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?        xxxxxx�?�?vb'vb'�?;�;��?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?      �?        9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?333333�?�������?              �?      �?              �?              �?      �?�Kh/��?�Kh/���?#>�Tr^�?���VC�?              �?������??4և���?L�Ϻ��?�g�`�|�?o0E>��?#�u�)��?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?�;�;�?�؉�؉�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?      �?              �?                      �?      �?      �?              �?      �?        �g�`�|�?o0E>��?9��8���?�q�q�?      �?      �?333333�?�������?      �?      �?              �?      �?              �?              �?              �?        n۶m۶�?%I�$I��?              �?=��<���?�a�a�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?              �?      �?        DDDDDD�?�����ݽ?�������?UUUUUU�?���Q��?{�G�z�?      �?      �?      �?        �������?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        �������?�������?wwwwww�?�?]t�E]�?F]t�E�?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�G         r                     @�����?�           8�@                                   �?yÏP�?�            �t@                                03�<@@+K&:~�?[             c@                                   �?Xny��?(            �N@                                 �H@>A�F<�?             C@                                  �?�t����?             A@                                 @B@�nkK�?             7@       ������������������������       �                     2@        	       
                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���!pc�?             &@        ������������������������       �                     �?                                  �;@�z�G��?             $@                                  �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                      @                                  �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �        3            �V@               =                    �?:���١�?p             f@               8                     �?�[�IJ�?            �G@              5                    �?      �?             C@                                ��";@��>4և�?             <@        ������������������������       �                      @        !       4                 �̾w@$��m��?             :@       "       '                 �|Y<@`�Q��?             9@        #       &                    �?      �?              @       $       %                  �}S@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        (       3                    �?@�0�!��?             1@       )       2                 p�i@@�θ�?	             *@       *       /                   �A@և���X�?             @       +       ,                 ���<@      �?             @        ������������������������       �                      @        -       .                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        6       7                 ��>Y@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        9       :                    �?�����H�?             "@       ������������������������       �                     @        ;       <                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        >       m                    �?
�e4���?Q             `@       ?       Z                     �?d�X^_�?I            �\@        @       O                    B@H.�!���?!             I@        A       N                 `f�D@�LQ�1	�?             7@       B       C                 ��I*@��S���?
             .@        ������������������������       �                     @        D       E                   �<@z�G�z�?             $@        ������������������������       �                     @        F       M                   @>@����X�?             @       G       L                 �|�?@���Q��?             @       H       I                 �|Y=@�q�q�?             @        ������������������������       �                     �?        J       K                 `fF<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        P       Y                 ���[@�����H�?             ;@       Q       X                    �?$�q-�?             :@       R       W                 `f�;@�C��2(�?             6@       S       V                   �K@r�q��?             (@        T       U                 ��:@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     �?        [       l                    �?P�2E��?(            @P@       \       k                   �*@�X�<ݺ?              K@       ]       ^                   �(@$�q-�?            �C@        ������������������������       �        	             ,@        _       `                 �|�<@H%u��?             9@        ������������������������       �                     "@        a       b                 �|�=@     ��?             0@        ������������������������       �                     �?        c       j                   �F@�r����?
             .@       d       i                   @D@z�G�z�?             $@       e       f                    @@�����H�?             "@        ������������������������       �                     @        g       h                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     &@        n       o                    :@X�Cc�?             ,@        ������������������������       �                     @        p       q                    5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        s                          @l���`��?�            �w@       t       �                    �?B�>�;Q�?�            �w@       u       �                    �?C؇eY�?�            �p@        v                        P��@�ucQ?-�?3            @U@        w       ~                 ���@      �?             8@       x       y                 03S@z�G�z�?
             .@        ������������������������       �                     �?        z       {                   �7@d}h���?	             ,@        ������������������������       �                      @        |       }                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     "@        �       �                    �?��7��?#            �N@       �       �                 �|Y=@\X��t�?             G@        �       �                    �?     ��?	             0@        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             (@       ������������������������       �                      @        �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�������?             >@        ������������������������       �                     @        �       �                 @a'@8����?             7@       �       �                 `�j@�q�q�?             5@       �       �                 X��A@�z�G��?             4@       �       �                 �;@�����?             3@       �       �                 03@�q�q�?             2@       �       �                 ��@�t����?             1@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@������?	             .@        ������������������������       �                     �?        �       �                    �?����X�?             ,@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�G�z�?             .@        �       �                    &@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���&@؇���X�?             @        ������������������������       �                     @        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �0@X��Oԣ�?t            @g@        ������������������������       �                     @        �       �                    �?�8��8��?o            �f@        �       �                 ���@�q�q�?
             .@        ������������������������       �                     �?        �       �                 �|�;@����X�?	             ,@       �       �                   �9@���|���?             &@       �       �                    8@�<ݚ�?             "@       �       �                   �6@����X�?             @       �       �                  �#@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@�FVQ&�?e            �d@        �       �                 �|Y=@`<)�+�?1            @S@       �       �                   �8@p���?             I@       �       �                   �7@ ��WV�?             :@       ������������������������       �                     7@        �       �                 `fF@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                 �|Y>@�>����?             ;@        �       �                  sW@�t����?
             1@        �       �                 ��,@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     &@        ������������������������       �        
             $@        �       �                   �3@`���i��?4             V@        �       �                   �1@�θ�?             *@        ������������������������       �                      @        �       �                 `�8"@���!pc�?             &@       �       �                   �2@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                   �:@Х-��ٹ?-            �R@        ������������������������       �                     <@        �       �                   �;@dP-���?             �G@        ������������������������       �                     �?        �       �                 @3�@���.�6�?             G@        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��) @ �#�Ѵ�?            �E@        ������������������������       �                     7@        �       �                 �|�>@ףp=
�?             4@       �       �                 pf� @r�q��?
             (@        ������������������������       �                     �?        �       �                    (@�C��2(�?	             &@        �       �                 �|Y=@z�G�z�?             @        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                          �?������?L             [@       �       �                    �?�BE����?)             O@        �       �                    �?      �?             $@       �       �                    �?X�<ݚ�?             "@       �       �                  S�-@����X�?             @        �       �                 03�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�	j*D�?!             J@       �       �                   �3@�P�*�?             ?@        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             ;@        ������������������������       �                     *@        �       �                 03�1@X�Cc�?             ,@        �       �                 ���.@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �                          �?؇���X�?             5@       �                          �?�KM�]�?             3@       �                        ��y'@�8��8��?	             (@        �       �                 P�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 $@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?*
;&���?#             G@        	                      ��*4@��<b���?             7@        
                        �1@      �?             @        ������������������������       �                      @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @�KM�]�?             3@                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@                                 �?���}<S�?             7@       ������������������������       �                     *@                                 @z�G�z�?             $@                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  �����?��܍��?Q��+Q�?W�v%jW�?Cy�5��?l(�����?�}�K�`�?C��6�S�?Cy�5��?������?�?<<<<<<�?d!Y�B�?�Mozӛ�?              �?�������?�������?      �?                      �?t�E]t�?F]t�E�?              �?333333�?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?              �?      �?      �?              �?      �?              �?      �?                      �?              �?/�袋.�?F]t�E�?���
b�?m�w6�;�?      �?      �?۶m۶m�?I�$I�$�?              �?�N��N��?vb'vb'�?��(\���?{�G�z�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?ZZZZZZ�?�������?ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?�������?�������?              �?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        ���-iK�?�%mI[��?�s���?�aܯK*�?�(\����?)\���(�?Nozӛ��?d!Y�B�?�������?�?      �?        �������?�������?              �?�$I�$I�?�m۶m��?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?              �?      �?        �q�q�?�q�q�?�؉�؉�?;�;��?]t�E�?F]t�E�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?                      �?_�^��?z�z��?��8��8�?�q�q�?�؉�؉�?;�;��?      �?        )\���(�?���Q��?      �?              �?      �?              �?�������?�?�������?�������?�q�q�?�q�q�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?              �?      �?        ��\��?��]�һ�?
�ZN��?���nT�?%��J?s�?m�}�3�?666666�?�������?      �?      �?�������?�������?      �?        I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        &C��6��?�y��!�?!Y�B�?��Moz��?      �?      �?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?�������?�������?      �?        d!Y�B�?8��Moz�?UUUUUU�?UUUUUU�?ffffff�?333333�?Q^Cy��?^Cy�5�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?        wwwwww�?�?      �?        �m۶m��?�$I�$I�?              �?      �?                      �?      �?              �?                      �?      �?        �������?�������?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        c�1�c�?�s�9�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?�m۶m��?�$I�$I�?]t�E]�?F]t�E�?9��8���?�q�q�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        >����?|���?S{����?��O���?\���(\�?{�G�z�?O��N���?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �Kh/��?h/�����?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        t�E]t�?]t�E]�?ى�؉��?�؉�؉�?      �?        F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        K~��K�?O贁N�?      �?        �����F�?W�+�ɵ?              �?���7���?Y�B��?UUUUUU�?UUUUUU�?              �?      �?        �/����?�}A_Ч?      �?        �������?�������?�������?UUUUUU�?              �?]t�E�?F]t�E�?�������?�������?      �?      �?      �?                      �?      �?              �?              �?        B{	�%��?{	�%���?)��RJ)�?���Zk��?      �?      �?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        vb'vb'�?;�;��?�RJ)���?�Zk����?              �?UUUUUU�?UUUUUU�?      �?        �m۶m��?%I�$I��?�������?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�k(���?(�����?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?      �?              �?      �?        ���,d!�?8��Moz�?��,d!�?��Moz��?      �?      �?              �?      �?      �?      �?                      �?�k(���?(�����?UUUUUU�?UUUUUU�?      �?                      �?      �?        ӛ���7�?d!Y�B�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�G         �                     @e�L��?�           8�@               Y                     �?x@����?�            �u@               P                   �J@���(�_�?k            �e@                               `V�9@�ӭ�a�?Y             b@        ������������������������       �                     @                                  �7@�:���?T             a@        ������������������������       �                     3@               %                   �?@�k��(A�?I            �]@        	                         x;K@Fx$(�?             I@       
                          �<@|��?���?             ;@        ������������������������       �                      @                                  �>@�����?             3@                               �|Y=@���Q��?	             .@        ������������������������       �                      @                                  �<@��
ц��?             *@        ������������������������       �                     @                                  @D@���Q��?             $@        ������������������������       �                     @                                  �I@z�G�z�?             @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               "                    �?��+7��?             7@                                  �?�t����?             1@       ������������������������       �                     (@                                `f�N@���Q��?             @        ������������������������       �                      @               !                    �?�q�q�?             @                                 �}S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        #       $                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        &       E                 x5Q@�M���?*             Q@       '       D                 0��M@ҳ�wY;�?             A@       (       1                 ���;@¦	^_�?             ?@        )       *                 03k:@8�Z$���?             *@        ������������������������       �                     @        +       ,                    �?z�G�z�?             $@        ������������������������       �                     �?        -       .                   �C@�<ݚ�?             "@        ������������������������       �                     @        /       0                    H@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        2       5                    �?b�2�tk�?             2@        3       4                 ��A@      �?              @        ������������������������       �                      @        ������������������������       �                     @        6       ;                    �?      �?             $@        7       :                    �?      �?             @       8       9                    C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        <       =                   �C@      �?             @        ������������������������       �                     �?        >       A                    �?���Q��?             @        ?       @                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       C                 �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       G                    �?l��\��?             A@       ������������������������       �        
             0@        H       I                    �?r�q��?	             2@        ������������������������       �                      @        J       O                    �?�z�G��?             $@       K       N                 Ј�U@      �?              @        L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                 �U'Q@ܷ��?��?             =@       ������������������������       �                     6@        S       T                    �?և���X�?             @        ������������������������       �                      @        U       V                   �K@z�G�z�?             @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �1@և���X�?k            �e@        [       \                    �?�}�+r��?             3@       ������������������������       �                     ,@        ]       ^                    #@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �                    L@����3��?_            �c@       a       |                    �?Fx$(�?Y            �b@        b       {                    :@��ϭ�*�?'             M@       c       d                    �?�����H�?            �F@        ������������������������       �                     @        e       z                    �?,���i�?            �D@       f       s                    �?6YE�t�?            �@@       g       j                   �9@�C��2(�?             6@        h       i                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �'@�}�+r��?             3@        ������������������������       �                     @        m       r                   �,@�8��8��?             (@       n       o                    B@�����H�?             "@       ������������������������       �                     @        p       q                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       y                   �E@���!pc�?             &@       u       x                   �;@�����H�?             "@        v       w                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        }       ~                 �|Y=@�nkK�?2             W@        ������������������������       �                     A@               �                   �*@ 	��p�?!             M@       �       �                    �?(N:!���?            �A@        ������������������������       �                     @        �       �                 �|�=@      �?             @@        �       �                    @�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   @D@�nkK�?             7@       ������������������������       �                     &@        �       �                 `f�)@�8��8��?             (@        ������������������������       �                      @        �       �                   �F@ףp=
�?             $@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     @        �       �                    @��,?S�?�            �v@        �       �                    @$��m��?             :@        ������������������������       �                     &@        �       �                    @���Q��?             .@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                      @        �       �                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�B���?�            u@        �       �                   @C@     ��?=             X@       �       �                    �?V�K/��?5            �S@        �       �                    �?���B���?             :@       �       �                    �?P���Q�?             4@        �       �                 ���,@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                 `�@1@�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @A@Fmq��?             �J@       �       �                   @1@���Q �?            �H@       �       �                    �?)O���?             B@       �       �                   �5@8�A�0��?             6@        �       �                   �3@؇���X�?             @       �       �                   !@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@��S���?             .@       �       �                 ��&@�n_Y�K�?
             *@       �       �                    ;@���!pc�?             &@       �       �                 03�!@և���X�?             @       �       �                   �7@      �?             @        ������������������������       �                      @        �       �                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?����X�?             ,@       �       �                    �?�θ�?             *@       �       �                 ���)@�q�q�?             "@        ������������������������       �                     @        �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @        ������������������������       �                     1@        �                          �?P�_��I�?�             n@       �       �                    �?      �?�             l@        �       �                 �=/@�<ݚ�?$             K@       �       �                   �7@@�0�!��?"            �I@        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��0{9�?            �G@        �       �                    �?�X�<ݺ?             2@       �       �                 �|Y?@��S�ۿ?             .@       �       �                 �|Y;@�����H�?             "@        ������������������������       �                     �?        �       �                 ���@      �?              @        ������������������������       �                     @        �       �                 p&�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                  ��@V�a�� �?             =@        ������������������������       �                     @        �       �                    �?���!pc�?             6@       �       �                 X��A@����X�?             5@       �       �                   @'@ҳ�wY;�?	             1@       ������������������������       �      �?             0@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �0@��O���?q            @e@        �       �                 pf�@      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �                 pFD!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �                         @@@���C"��?l            �d@       �                          �? �	.��?V            ``@       �                       �!&B@�|K��2�?U             `@       �                       �|�=@�[|x��?S            �_@       �                       �|Y=@@-�_ .�?K            �[@       �                          �?�F��O�?7            @R@       �       �                   �:@�U�=���?1            �P@       �       �                 @3�@@9G��?'            �H@       ������������������������       �                     :@        �       �                 0S5 @���}<S�?             7@        �       �                   �2@      �?              @        ������������������������       �                     �?        �       �                   �3@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     .@                               pf� @@�0�!��?
             1@       ������������������������       �                     "@                              ���)@      �?              @                               �;@      �?             @        ������������������������       �                      @                                �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        	                         5@؇���X�?             @        
                      �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@                                �?@������?             .@                                �>@      �?              @                              (Se!@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                              pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?؇���X�?             @                             ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �        	             1@        �t�b�+z      h�h)h,K ��h.��R�(KMKK��h^�B�  v�S(��?��X��?�f��o��?�L�Ȥ�?�wK�?��?DZ/`��?��8��8�?9��8���?      �?        �8R4��?C�q���?              �?~ylE�p�?A�Iݗ��?R���Q�?ףp=
��?	�%����?{	�%���?              �?Q^Cy��?^Cy�5�?333333�?�������?      �?        �;�;�?�؉�؉�?      �?        �������?333333�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        Y�B��?zӛ����?�?<<<<<<�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?<<<<<<�?�������?�������?�������?�RJ)���?��Zk���?;�;��?;�;��?              �?�������?�������?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?      �?              �?9��8���?�8��8��?      �?      �?      �?                      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?        �������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?------�?              �?UUUUUU�?�������?              �?333333�?ffffff�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��=���?a���{�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?(�����?�5��P�?              �?�������?�������?              �?      �?        ��N��N�?'vb'vb�?ףp=
��?R���Q�?|a���?����=�?�q�q�?�q�q�?              �?8��18�?�����?e�M6�d�?'�l��&�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?(�����?�5��P�?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?t�E]t�?F]t�E�?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?                      �?              �?�Mozӛ�?d!Y�B�?      �?        ������?�{a���?|�W|�W�?�A�A�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?              �?        �ˠT�?����|��?vb'vb'�?�N��N��?              �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?W.��eZ�?�F��h��?      �?      �?�Z܄��?�ґ=�?ى�؉��?��؉���?�������?ffffff�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�x+�R�?~�	�[�?9/����?����>4�?9��8���?��8��8�?/�袋.�?颋.���?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�?�������?;�;��?ى�؉��?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?                      �?              �?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?      �?                      �?      �?        |;H|;H�?$�$��?      �?      �?9��8���?�q�q�?ZZZZZZ�?�������?      �?      �?              �?      �?        m�w6�;�?L� &W�?��8��8�?�q�q�?�������?�?�q�q�?�q�q�?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        ��{a�?a���{�?      �?        F]t�E�?t�E]t�?�m۶m��?�$I�$I�?�������?�������?      �?      �?      �?              �?              �?                      �?�������?�?      �?      �?      �?        �������?333333�?      �?      �?              �?      �?                      �?w%jW�v�?KԮD�J�?@u���?�U���g�?2g�s��?sƜ1g̹?]�u]�u�?EQEQ�?S�n0E�?к����?�իW�^�?�P�B�
�?�M6�d��?e�M6�d�?������?9/���?      �?        ӛ���7�?d!Y�B�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        ZZZZZZ�?�������?      �?              �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        wwwwww�?�?      �?      �?333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?      �?      �?              �?                      �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMIhvh)h,K ��h.��R�(KMI��h}�B@R         N                    �?�t����?�           8�@                                   �?�9��L~�?^            �b@                                `�@1@�C��2(�?)            �P@                                   �?�E��ӭ�?             2@                                  �?�8��8��?             (@       ������������������������       �                     @                                P��+@z�G�z�?             @        ������������������������       �                      @        	       
                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�q�q�?             @                               �&�)@���Q��?             @        ������������������������       �                     �?                                  �-@      �?             @        ������������������������       �                      @                                ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                  �H@@��8��?             H@       ������������������������       �                     D@                                   �?      �?              @                                   �?      �?             @                               ,w�U@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               -                 pF�#@�t����?5            @U@               "                   �5@�#-���?            �A@                !                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       $                 ���@�FVQ&�?            �@@        ������������������������       �                     ,@        %       (                 �|Y=@�KM�]�?             3@        &       '                   @@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        )       ,                   @@��S�ۿ?
             .@        *       +                 �|�=@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     $@        .       I                     @� �	��?             I@       /       D                     �?�D����?             E@       0       C                   �H@X�<ݚ�?             B@       1       2                 �|Y<@���!pc�?             6@        ������������������������       �                     @        3       >                    �?ҳ�wY;�?             1@       4       ;                 `f�A@�q�q�?             (@       5       :                 X�,@@      �?              @       6       7                 �ܵ<@���Q��?             @        ������������������������       �                     �?        8       9                 ��2>@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        <       =                 @�Cq@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       @                   @H@z�G�z�?             @        ������������������������       �                     �?        A       B                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        E       F                 ���@@r�q��?             @       ������������������������       �                     @        G       H                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        J       M                    �?      �?              @        K       L                   �3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       �                   �3@�钹H��?^           ��@        P       �                    @��o	��?D             ]@       Q       v                    �?8�$�>�?4            �U@       R       S                    �?
;&����?             G@        ������������������������       �                     @        T       q                    6@�G��l��?             E@       U       n                    �?���Q��?            �A@       V       ]                    �?J�8���?             =@        W       X                   �1@z�G�z�?             @        ������������������������       �                     �?        Y       \                 ��!@      �?             @       Z       [                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ^       a                     @      �?             8@        _       `                   �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        b       g                   �1@���y4F�?             3@        c       f                   �0@      �?              @        d       e                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        h       m                 0S5 @���!pc�?             &@        i       j                   �2@      �?             @        ������������������������       �                      @        k       l                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       p                   �2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        r       s                     �?؇���X�?             @        ������������������������       �                     �?        t       u                   �1@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        w       ~                    �?z�G�z�?             D@        x       y                     @�t����?             1@       ������������������������       �                     $@        z       {                    �?����X�?             @        ������������������������       �                     @        |       }                 `f7@      �?             @       ������������������������       �                      @        ������������������������       �                      @               �                    )@��+7��?             7@       �       �                    �?�KM�]�?             3@       ������������������������       �                     *@        �       �                    �?�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             >@        �       �                    @ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    *@��
ц��?             *@       �       �                    @�z�G��?             $@        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                     @�/e�U��?           �{@        �       �                    �?      �?v             g@       �       �                    �?*��w\��?\            �b@        �       �                    :@=QcG��?            �G@        �       �                   �3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �B@�Ń��̧?             E@       ������������������������       �                     9@        �       �                   @C@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    �?��[�8��?B            �Y@        ������������������������       �                     �?        �       �                     �?�C+����?A            @Y@       �       �                    �?���Q �?!            �H@       �       �                   �B@�z�G��?             D@       �       �                   �A@���Q��?             >@       �       �                   �>@�q�q�?             ;@       �       �                   @>@և���X�?             5@       �       �                 �̌*@�q�q�?             2@        ������������������������       �                     @        �       �                 `fF<@և���X�?
             ,@       �       �                   @L@�eP*L��?             &@       �       �                    H@      �?              @       �       �                 �|�<@      �?             @        ������������������������       �                     �?        �       �                 �|�?@���Q��?             @        ������������������������       �                     �?        �       �                   �C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    =@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��<R@      �?              @       �       �                   �C@z�G�z�?             @        ������������������������       �                      @        �       �                  x#J@�q�q�?             @        ������������������������       �                     �?        �       �                 �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ,@4��?�?              J@       �       �                 `f�)@�חF�P�?             ?@        ������������������������       �        	             (@        �       �                   �A@�d�����?             3@        �       �                 �|Y<@      �?              @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        �       �                    @@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        �       �                   �F@�C��2(�?             &@       �       �                   @D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     5@        �       �                   �M@��R[s�?            �A@       �       �                    F@     ��?             @@       �       �                    B@�+e�X�?             9@       �       �                    �?R���Q�?             4@       ������������������������       �                     1@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                          �?�����D�?�            @p@        �                          �?�ʻ����?.             Q@       �       �                 ��@�~8�e�?$            �I@        �       �                    �?@�0�!��?             1@       �       �                 ���@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 pff@����X�?             @       �       �                 �|�9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�ʻ����?             A@        ������������������������       �                     @        �                         �>@d��0u��?             >@       �       �                 ��&@l��
I��?             ;@       �       �                   �@�r����?
             .@        �       �                 �&B@      �?             @       �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �                          4@      �?             (@       �       �                   �:@      �?              @        ������������������������       �                     �?        �                           �?؇���X�?             @        ������������������������       �                     @                                �.@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              �|�:@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        	      D                ���5@     ��?v             h@       
      ?                   �?�L���?r             g@             6                ���"@d#,����?e            �d@                                �?@�+9\J�?Z            �b@                              �|Y=@؇���X�?             5@                               ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              X�I@�KM�]�?             3@                             ���@�t����?             1@        ������������������������       �                      @                              ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @                                �7@����?K            @`@        ������������������������       �                    �A@                              ���@<����?7            �W@        ������������������������       �        	             2@                                @8@�s�c���?.            @S@                              03@      �?             @        ������������������������       �                      @        ������������������������       �                      @               1                @3�@�F��O�?,            @R@       !      "                �|Y=@X�EQ]N�?            �E@        ������������������������       �                     .@        #      0                  �C@�>4և��?             <@       $      %                pf�@�E��ӭ�?             2@        ������������������������       �                     @        &      /                   B@�q�q�?
             (@       '      .                  @@@���|���?	             &@       (      )                  �@���Q��?             $@        ������������������������       �                     @        *      +                �|�>@؇���X�?             @        ������������������������       �                     @        ,      -                �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        2      5                �|Y<@(;L]n�?             >@        3      4                  �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        7      <                �|�=@d}h���?             ,@       8      9                  �<@�C��2(�?	             &@       ������������������������       �                     @        :      ;                �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =      >                  �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @      C                pf� @P���Q�?             4@        A      B                ��Y@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        E      H                   �?և���X�?             @        F      G                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMIKK��h^�B�  G�+J>�?r%�k���?��o�7��?��d�?F]t�E�?]t�E�?r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?      �?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�������?�������?�A�A�?_�_�?      �?      �?      �?                      �?>����?|���?      �?        �k(���?(�����?      �?      �?      �?                      �?�������?�?�������?�������?      �?      �?      �?              �?        �Q����?)\���(�?�0�0�?z��y���?r�q��?�q�q�?t�E]t�?F]t�E�?              �?�������?�������?�������?�������?      �?      �?�������?333333�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?                      �?�������?�������?              �?      �?      �?              �?      �?              �?        �������?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?333333�?�������?              �?      �?                      �?PuPu�?_�_��?������?���{�?�5eMYS�?6eMYS��?�Mozӛ�?Y�B��?              �?1�0��?��y��y�?333333�?�������?�rO#,��?|a���?�������?�������?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?333333�?�������?      �?                      �?6��P^C�?(������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?�������?�������?�?<<<<<<�?              �?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?        Y�B��?zӛ����?(�����?�k(���?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?      �?              �?        �������?�������?�������?�������?      �?        �;�;�?�؉�؉�?ffffff�?333333�?      �?      �?      �?                      �?      �?                      �?      �?        �^����?�B�I .�?      �?      �?l}0T��?(ɟWY�?AL� &W�?x6�;��?�������?333333�?      �?                      �?�a�a�?��<��<�?              �?�?�?      �?                      �?�?�������?      �?        &���?��g����?9/����?����>4�?ffffff�?333333�?333333�?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?t�E]t�?]t�E�?      �?      �?      �?      �?              �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        �q�q�?r�q��?              �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�N��N��?ى�؉��?�Zk����?��RJ)��?      �?        Cy�5��?y�5���?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?      �?              �?      �?]t�E�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?        PuPu�?X|�W|��?      �?      �?���Q��?R���Q�?333333�?333333�?              �?      �?        333333�?�������?              �?      �?                      �?      �?        z�z��?z�z��?�������?<<<<<<�?�������?222222�?�������?ZZZZZZ�?�������?�������?      �?                      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�������?<<<<<<�?              �?DDDDDD�?wwwwww�?Lh/����?h/�����?�������?�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?                      �?�?�?              �?      �?              �?      �?}���g�?L�Ϻ��?I����H�?��[���?�vV;��?��JL%��?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?�k(���?(�����?<<<<<<�?�?      �?        9��8���?�q�q�?      �?      �?      �?              �?        ~�~��? �����?      �?        ���%N�?�X�0Ҏ�?      �?        �����?�cj`?      �?      �?              �?      �?        �իW�^�?�P�B�
�?w�qG�?qG�wĽ?      �?        �$I�$I�?�m۶m��?�q�q�?r�q��?      �?        �������?�������?]t�E]�?F]t�E�?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?        I�$I�$�?۶m۶m�?]t�E�?F]t�E�?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ffffff�?�������?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?        �t�bubhhubehhub.